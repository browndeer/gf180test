* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_39_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3691__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout56_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5968__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4640__B2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6845_ _0072_ net207 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6776_ _0406_ net165 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4243__I1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ mod.registers.r4\[12\] _0974_ _0980_ mod.registers.r14\[12\] _1016_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ _2503_ _2561_ _2563_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4943__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _2479_ _2515_ _2520_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4609_ _1126_ _1315_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5589_ _2115_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5120__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6629__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6335__I _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6779__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A3 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4934__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3627__C _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3370__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5111__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4870__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4870__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _1899_ _1977_ _1980_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_91_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__I1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ _0912_ _0913_ _0914_ _0915_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4891_ _1848_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6630_ _0263_ net83 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3842_ _0714_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ _0194_ net56 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3773_ mod.registers.r11\[8\] _0799_ _0800_ mod.registers.r6\[8\] _0801_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4925__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5512_ mod.registers.r7\[3\] _2418_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6492_ _0125_ net117 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5443_ _2333_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _2304_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5350__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__C1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3361__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4325_ _1046_ _1038_ _1351_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3361__B2 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout105 net109 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout127 net129 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout138 net139 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4256_ _1177_ _3129_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5102__A2 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ _1175_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4613__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _0055_ net191 mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3719__A3 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _0389_ net180 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4472__S0 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3655__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4852__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4907__A2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__B _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ _1130_ _1137_ _0735_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5090_ _1794_ _2082_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4041_ _1064_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3646__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _2707_ _2750_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5399__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _1899_ _1960_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4071__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4874_ _3099_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6613_ _0246_ net46 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3825_ _0844_ _0847_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _0177_ net98 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3756_ _3139_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3582__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3582__B2 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _3085_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3687_ _0714_ _0710_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ mod.registers.r5\[8\] _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3334__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ mod.registers.r4\[5\] _2311_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3885__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _1080_ _1009_ _1024_ _1246_ _1335_ _1234_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ mod.registers.r2\[14\] _2264_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5087__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4239_ _1037_ _1196_ _0643_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_28_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4834__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3637__A2 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5938__B _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4062__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A4 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6339__B2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5229__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3573__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__A2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5899__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6497__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5002__A1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3610_ mod.registers.r13\[2\] _3140_ _3144_ mod.registers.r1\[2\] _0637_ _0638_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4590_ _1598_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5553__A2 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3564__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _0436_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _2892_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3472_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5305__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5211_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6191_ _2903_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ mod.registers.r1\[4\] _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3619__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4024_ _1049_ _1050_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__I _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__B _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _2721_ _2729_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6433__I _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4926_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _0622_ _1880_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ _0793_ _0795_ _0798_ _0801_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__A3 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _1804_ _1814_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6527_ _0160_ net88 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4752__B1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__I _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3739_ _0623_ _0625_ _0627_ _0629_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4752__C2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ mod.des.des_dout\[24\] net9 _3071_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5409_ _2346_ _2347_ _2349_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6389_ _2270_ _2567_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3858__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5480__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3491__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5783__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3794__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3794__B2 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3546__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5422__I _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout173_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__S _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3482__B1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__B _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5760_ mod.registers.r12\[8\] _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5774__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4711_ _3105_ _1726_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _2270_ _2442_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4642_ _1653_ _1658_ _1659_ _1662_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_30_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5526__A2 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3537__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I0 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4573_ _1518_ _1447_ _1389_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _1802_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3524_ mod.registers.r1\[4\] _0483_ _0551_ mod.registers.r7\[4\] _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6243_ _1133_ _2658_ _2937_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3455_ _3230_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout86_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6174_ _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6512__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3386_ mod.instr_2\[16\] _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3561__B _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ mod.des.des_dout\[23\] _2105_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ mod.pc0\[13\] _1889_ _1961_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _0902_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5958_ _2721_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5765__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _1736_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5889_ _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3528__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3528__B2 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4411__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4567__B _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3464__B1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3464__C2 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__B2 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5508__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6535__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3240_ _3096_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6248__I _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5444__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _0088_ net102 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3470__A3 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5812_ _2598_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _0019_ net158 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5743_ _2477_ _2570_ _2574_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4940__B mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _2493_ _2528_ _2530_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4625_ _1405_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6172__A2 _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4231__I _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _1278_ _1480_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3507_ mod.registers.r6\[5\] _0417_ _3226_ mod.registers.r2\[5\] _3230_ mod.registers.r1\[5\]
+ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _1506_ _1510_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _2890_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3438_ mod.registers.r4\[6\] _3177_ _3181_ mod.registers.r2\[6\] _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4486__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A1 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6158__I _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6157_ net13 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _3200_ _3202_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3694__B1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _2101_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6088_ _2825_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ mod.pc\[12\] _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A1 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3997__B2 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3749__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__B _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4410__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4174__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3921__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput20 net20 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5674__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__I _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_223 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_234 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_245 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5426__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_256 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_267 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_278 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3437__B1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_289 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3988__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3988__B2 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4316__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout136_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6154__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _0567_ _0588_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5390_ mod.registers.r5\[0\] _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5901__A2 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ _1263_ _1368_ _1267_ _1234_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4986__I mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _1290_ _1298_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5665__A1 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _2767_ _2766_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5417__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4654__C _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3979__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _0071_ net211 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6700__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__B _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ _0405_ net167 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3987_ mod.registers.r9\[12\] _0977_ _0522_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5726_ mod.registers.r11\[12\] _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5657_ mod.registers.r10\[2\] _2517_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6850__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ _1405_ _1632_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5588_ _2385_ _2464_ _2469_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4539_ _1130_ _1313_ _1217_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5656__A1 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _2889_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4845__B _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5408__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3975__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4395__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5895__A1 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3416__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3370__A2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6447__I0 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__A2 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6723__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__I2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3910_ _0922_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _1653_ _1607_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3841_ _0445_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3772_ _0464_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6560_ _0193_ net94 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5511_ _2340_ _2416_ _2421_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6491_ _0124_ net115 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4138__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5442_ _2331_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5886__A1 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ _2302_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3897__B1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3897__C2 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4324_ _0945_ _0956_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3361__A2 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout106 net109 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout117 net118 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4255_ _1214_ _1227_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xfanout139 net140 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4186_ _1182_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A1 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5810__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6372__S _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__B1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _0054_ net191 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3795__I _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ _0388_ net155 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4472__S1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5709_ _2487_ _2549_ _2552_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6118__A2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6689_ _0322_ net54 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5515__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4559__C _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5629__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3591__A2 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__I _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__B2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4040_ _1065_ _1066_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3646__A3 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4056__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5991_ _2710_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ mod.pc0\[6\] _1909_ _1961_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_33_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _0000_ _0675_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6348__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4359__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6612_ _0245_ net51 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3824_ _0848_ _0849_ _0850_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3755_ mod.registers.r9\[8\] _0781_ _0782_ mod.registers.r3\[8\] _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6543_ _0176_ net100 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6619__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3582__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ mod.des.des_dout\[30\] net2 _3084_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3686_ _3134_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5859__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2333_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3334__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5356_ _2145_ _2310_ _2312_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _1264_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _2225_ _2263_ _2266_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4238_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4169_ _0834_ _1109_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4350__S _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4522__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6275__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__S0 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4038__B1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A3 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5002__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3540_ mod.pc_2\[4\] _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3564__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4761__A1 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3471_ _3166_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5210_ mod.des.des_dout\[32\] _2187_ _2205_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6190_ _2890_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _2117_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ mod.ins_ldr_3 mod.valid_out3 net15 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4816__A2 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4023_ mod.registers.r4\[14\] _0974_ _0975_ mod.registers.r11\[14\] _1051_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3403__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _1926_ _2735_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4925_ _0532_ _0536_ _3092_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ _1735_ _1863_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3807_ _0783_ _0785_ _0787_ _0789_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4787_ mod.ldr_hzd\[13\] _1795_ _1803_ mod.ldr_hzd\[12\] _1799_ mod.ldr_hzd\[15\]
+ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6526_ _0159_ net94 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4752__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3738_ mod.pc_2\[2\] _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4752__B2 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ _3074_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3669_ mod.registers.r12\[1\] _0694_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5408_ mod.registers.r5\[4\] _2348_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6388_ _3032_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5339_ _2097_ _2269_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6257__A1 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4268__B1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5014__B _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5480__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3491__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3491__B2 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5232__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3794__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3546__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout166_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5223__A2 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4054__I _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _1728_ _1733_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ _2511_ _2534_ _2539_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4641_ _1469_ _1666_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3537__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__A1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _1518_ _1447_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6311_ _1755_ _2974_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3523_ _0430_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6242_ mod.pc_1\[0\] _2936_ _2822_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3454_ mod.registers.r13\[6\] _0480_ _0481_ mod.registers.r14\[6\] _0482_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ mod.valid1 _2653_ _2661_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3385_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6239__A1 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _2129_ _1877_ _2122_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout79_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ _2069_ _1868_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4006_ _0829_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6411__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _2720_ _1856_ _1739_ _1840_ _2715_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1876_ _1914_ _1916_ _1917_ _1931_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4973__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4839_ _1728_ _1859_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3528__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _0142_ net87 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__A1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3464__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3464__B2 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A2 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3767__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5433__I _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__S _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4493__B _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ _0087_ net103 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _2596_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6791_ _0018_ net159 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ mod.registers.r12\[1\] _2572_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ mod.registers.r10\[8\] _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5608__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4624_ _1635_ _1636_ _1639_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_129_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5380__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _1581_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3506_ mod.registers.r5\[5\] _0423_ _3219_ mod.registers.r4\[5\] _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4486_ _1511_ _1513_ _1281_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__B _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2923_ _2926_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3437_ mod.registers.r3\[6\] _3171_ _0464_ mod.registers.r6\[6\] _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6156_ mod.des.des_dout\[16\] _2872_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3368_ _3203_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__A1 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__B2 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _2662_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3299_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _1985_ _2047_ _2053_ _1843_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input11_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6174__I _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4246__I0 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4946__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3749__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5371__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3382__B1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3921__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 net21 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3685__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_224 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_235 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_246 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_257 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_268 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_279 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3437__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3437__B2 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3988__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6033__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5428__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout129_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ _1264_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_4_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4271_ _1297_ _0952_ _1296_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6259__I _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ mod.pc\[8\] _1993_ _1890_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input3_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5417__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3443__A4 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6843_ _0070_ net211 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4928__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _0404_ net167 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4928__B2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3986_ mod.registers.r6\[12\] _0960_ _0968_ mod.registers.r10\[12\] _1014_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3567__B _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5725_ _2543_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _2477_ _2515_ _2519_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _1121_ _1632_ _1634_ _1402_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5587_ mod.registers.r8\[15\] _2465_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4538_ _1379_ _1419_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3903__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5105__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ _1120_ _1488_ _1496_ _1401_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_89_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _2907_ _2915_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ mod.instr\[12\] _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__I _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6456__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6081__A2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4395__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6079__I _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5647__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6447__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4327__I _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4083__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4473__I3 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ _0804_ _0861_ _0867_ _0497_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__5583__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _3163_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5510_ mod.registers.r7\[2\] _2418_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _0123_ net118 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5335__A1 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5372_ _2209_ _2316_ _2321_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3897__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3897__B2 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4323_ _1041_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout107 net109 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout129 net137 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4254_ _1230_ _1255_ _1280_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _1186_ _1198_ _1203_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5621__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4237__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A2 _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3821__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3821__B2 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6826_ _0053_ net193 mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5574__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6757_ _0387_ net152 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5068__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3969_ _0806_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5708_ mod.registers.r11\[5\] _2550_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6688_ _0321_ net105 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6374__I0 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _2224_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3337__B1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4147__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3591__A3 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3879__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4540__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout196_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__I _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3500__B1 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4056__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5990_ _2748_ _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6840__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4056__B2 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4872_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6611_ _0244_ net52 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4359__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ mod.registers.r9\[9\] _0781_ _0516_ mod.registers.r12\[9\] _0851_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5556__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ _0175_ net98 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3754_ _3170_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6473_ _3077_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3685_ _3178_ _0710_ mod.registers.r1\[1\] _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5424_ _2331_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5355_ mod.registers.r4\[4\] _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3334__A3 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _1182_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4676__B _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5286_ mod.registers.r2\[13\] _2264_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4237_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4047__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4099_ _1010_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5795__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _0036_ net162 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4755__C1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A2 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6713__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4522__A2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3730__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6275__A2 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6863__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4381__S1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4038__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__B2 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4589__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__B1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3549__B1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4761__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4340__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout111_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout209_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3470_ _3199_ _0486_ _0496_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3721__B1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4496__B _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _2080_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4277__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ mod.registers.r14\[14\] _0980_ _0965_ mod.registers.r1\[14\] _1050_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ _1942_ _1943_ mod.pc\[4\] _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4924_ _1941_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4855_ _0730_ _0503_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _0507_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ mod.ldr_hzd\[14\] _1802_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6736__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _0158_ net88 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3737_ _0562_ _0608_ _0618_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__4752__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4250__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ mod.des.des_dout\[23\] net8 _3071_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3668_ _3232_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _2333_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5701__A1 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ mod.des.des_dout\[12\] net10 _3016_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6886__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3599_ mod.registers.r11\[2\] _0626_ _0571_ mod.registers.r2\[2\] _0627_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3712__B1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5338_ _2298_ _2089_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4268__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _2167_ _2251_ _2255_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3491__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3779__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6193__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3951__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6087__I _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__RN _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6609__CLK net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6420__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout159_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6759__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4640_ _1654_ _1315_ _1483_ _1279_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _1594_ _1595_ _1596_ _1185_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4734__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I2 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6310_ _2976_ _2980_ _2981_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3522_ mod.registers.r2\[4\] _0477_ _0488_ mod.registers.r9\[4\] mod.registers.r13\[4\]
+ _0480_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6241_ _2892_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3453_ _3212_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6172_ _2887_ _2826_ _2888_ _2828_ _2889_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3384_ mod.instr_2\[17\] _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_69_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _0766_ _2123_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5054_ mod.pc\[13\] _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4005_ _0986_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4245__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ mod.pc\[1\] _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_52_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _1899_ _1926_ _1930_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5887_ _2655_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4973__A2 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _1862_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _1793_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3933__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6508_ _0141_ net115 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _3064_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3324__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3464__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3621__C1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4716__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5714__I _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _2370_ _2610_ _2615_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6790_ _0017_ net158 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ _2470_ _2570_ _2573_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4955__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ _2516_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _1334_ _1642_ _1650_ _1281_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5904__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _0727_ _0762_ _0772_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3853__B _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3391__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ mod.registers.r7\[5\] _0431_ _3224_ mod.registers.r3\[5\] _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4485_ _1361_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _0695_ _2924_ _2920_ mod.instr\[14\] _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3436_ _3172_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6155_ mod.instr\[16\] _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ mod.instr_2\[14\] _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3694__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ mod.des.des_dout\[21\] _2105_ _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ mod.instr\[0\] _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3298_ _3146_ _3148_ _3133_ _3135_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_73_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5037_ _1985_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4643__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6396__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__A2 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4246__I1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4946__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6190__I _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__I _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3382__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3382__B2 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5534__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3921__A3 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3685__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_225 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4594__B _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_236 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_247 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_258 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_269 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4634__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3437__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__B _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5362__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4488__C _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _0952_ _1296_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6311__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6476__S _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4873__A1 _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6842_ _0069_ net212 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6773_ _0403_ net167 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4928__A2 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3985_ mod.registers.r11\[12\] _0975_ _0963_ mod.registers.r3\[12\] _1013_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5724_ _2541_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5655_ mod.registers.r10\[1\] _2517_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4606_ _1387_ _1633_ _1301_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5586_ _2382_ _2464_ _2468_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4537_ _1285_ _1435_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3903__A3 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5354__I _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6302__A1 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _1492_ _1495_ _1293_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6207_ _3119_ _2910_ _2913_ mod.instr\[8\] _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3419_ _0439_ _0444_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4399_ _1394_ _1403_ _1406_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ _2862_ _2863_ _2864_ _2855_ _2856_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6185__I _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6069_ mod.pc_1\[8\] _2812_ _2807_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3419__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5041__A1 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3658__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4855__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6095__I mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__C1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3512__I mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6028__C _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__A1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4083__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4343__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ mod.registers.r14\[8\] _0796_ _0797_ mod.registers.r10\[8\] _0798_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _2216_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6383__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__B _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5371_ mod.registers.r4\[11\] _2317_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _1007_ _1010_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4253_ _1177_ _3129_ _1176_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfanout119 net138 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4184_ _1211_ _1199_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6825_ _0052_ net193 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3968_ mod.registers.r5\[13\] _0559_ _0816_ mod.registers.r6\[13\] mod.registers.r14\[13\]
+ _0820_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6756_ _0386_ net187 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5707_ _2483_ _2549_ _2551_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6687_ _0320_ net94 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3899_ mod.registers.r6\[10\] _0816_ _0817_ mod.registers.r13\[10\] _0927_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5638_ _2503_ _2504_ _2506_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6374__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3337__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3337__B2 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5569_ _2444_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6642__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5014__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3576__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6792__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6365__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3879__A2 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3500__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3500__B2 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4056__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _1942_ _1943_ mod.pc\[6\] _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4871_ _1611_ _1628_ _1731_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6202__B1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _0243_ net53 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3822_ mod.registers.r4\[9\] _0628_ _0784_ mod.registers.r13\[9\] _0850_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5556__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _0174_ net100 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3753_ _3151_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4801__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _3083_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3684_ _0711_ _0635_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5118__B _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5354_ _2304_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6515__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4305_ _1297_ _1315_ _1321_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _2217_ _2263_ _2265_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4819__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4236_ _0747_ _0748_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _0562_ _0738_ _0746_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6665__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4098_ _1039_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5244__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__I _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _0035_ net162 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4755__B1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6739_ _0369_ net151 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3730__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5483__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__A1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A1 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__B2 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3549__A1 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3549__B2 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout90 net97 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6538__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout104_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5171__B1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3721__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3721__B2 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6688__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5070_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ mod.registers.r7\[14\] _0962_ _0960_ mod.registers.r6\[14\] _0959_ mod.registers.r13\[14\]
+ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__6484__S _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5226__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5777__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _2728_ _2706_ _2734_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4923_ mod.pc0\[5\] _1835_ _1845_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4017__B _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ _0447_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3805_ mod.pc_2\[8\] _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4785_ _1763_ _1802_ _1812_ _1781_ _1804_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3736_ _3199_ _0444_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6524_ _0157_ net116 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _3073_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3667_ _3220_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ _2331_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6386_ _3031_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3598_ _3163_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3712__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5337_ _2085_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3712__B2 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ mod.registers.r2\[6\] _2252_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4268__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4219_ _1246_ _1208_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _2177_ _2022_ _2196_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5217__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3779__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3779__B2 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__I0 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3951__B2 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3703__A1 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__B1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3520__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5447__I _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ _1453_ _1597_ _1456_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5931__A2 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I3 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ mod.registers.r10\[4\] _0547_ _0548_ mod.registers.r11\[4\] _0549_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _2930_ _2935_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ _3233_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6171_ _2649_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3383_ _3214_ _3227_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5122_ _2120_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ _2037_ _2066_ _2067_ _1868_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4004_ _1025_ _1026_ _1027_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_66_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5131__B _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _2705_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4422__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4906_ mod.pc0\[4\] _1887_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5886_ _2664_ _2666_ _2660_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _1735_ _1863_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4261__I _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6853__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3933__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6507_ _0140_ net119 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3933__B2 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3719_ _0645_ _0738_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4699_ _3109_ _1724_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ mod.des.des_dout\[15\] net18 _3061_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6369_ _3016_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5438__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5989__A2 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4110__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A1 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3621__B1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3621__C2 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6098__I mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4101__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout171_I net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5886__B _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6876__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ mod.registers.r12\[0\] _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5671_ _2514_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4622_ _1322_ _1643_ _1644_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5904__A2 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4553_ _1433_ _1435_ _1436_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3504_ _0528_ _0529_ _0530_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4484_ _1082_ _1231_ _1136_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5668__A1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3435_ _0458_ _0459_ _0461_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6223_ _2923_ _2925_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4030__B _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ _2874_ _2875_ _2876_ _2867_ _2868_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout84_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3366_ _3218_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _1133_ _2107_ _2109_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _2069_ _2819_ _2823_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3297_ _3147_ _3148_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5036_ mod.pc_2\[12\] _1074_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_100_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5840__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3851__B1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6396__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _1868_ _1928_ _2655_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5869_ _2652_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4159__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3906__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3382__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput23 net23 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3335__I _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3685__A3 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5550__I _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_226 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_237 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_248 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_259 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5831__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__I _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4873__A2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _0068_ net212 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4389__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6772_ _0402_ net168 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ mod.pc_2\[12\] _0834_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5050__A2 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ _2501_ _2555_ _2560_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5654_ _2470_ _2515_ _2518_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _1351_ _1162_ _1169_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5585_ mod.registers.r8\[14\] _2465_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4010__B1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5635__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4561__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ _0761_ _0734_ _0735_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _1432_ _1437_ _1494_ _1441_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6302__A2 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4313__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6206_ _2907_ _2914_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4313__B2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ mod.funct3\[2\] _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4398_ _1182_ _1418_ _1422_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ mod.des.des_dout\[11\] _2860_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3349_ mod.instr_2\[16\] _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A1 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _2804_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4616__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ mod.pc0\[11\] mod.pc\[11\] _1834_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4001__B1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4068__B1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__B1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout134_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5455__I _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _2202_ _2316_ _2320_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4321_ _1119_ _3130_ _1285_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ _1257_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xfanout109 net112 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4183_ _1205_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5190__I _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4059__B1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5271__A2 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout47_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6824_ _0051_ net182 mod.rd_3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ _0385_ net153 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3967_ _0989_ _0990_ _0993_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5706_ mod.registers.r11\[4\] _2550_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6686_ _0319_ net98 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ _0923_ _0924_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5637_ mod.registers.r9\[12\] _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4534__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3337__A2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5568_ _2357_ _2452_ _2457_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _1358_ _1543_ _1544_ _1236_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5499_ mod.registers.r6\[15\] _2409_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6196__I _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5014__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5984__B _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__B2 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3576__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4773__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3523__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3500__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4782__C _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__A1 _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ _1876_ _1877_ _1878_ _1852_ _1895_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_60_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6202__A1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6202__B2 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ mod.registers.r7\[9\] _0632_ _0788_ mod.registers.r15\[9\] _0849_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3567__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _0173_ net116 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3752_ _0500_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6471_ mod.des.des_dout\[29\] net19 _3079_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3683_ _3174_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5422_ _2183_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _2302_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _1322_ _1324_ _1328_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6010__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5284_ mod.registers.r2\[12\] _2264_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4235_ _0673_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4166_ _0645_ _0525_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4097_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4264__I _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _0034_ net162 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4999_ _1966_ _1999_ _2000_ _1997_ _2017_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6738_ _0368_ net151 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3802__I0 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _0302_ net105 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4213__B _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5095__I _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4507__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5180__A1 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5823__I _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3730__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__A2 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3797__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3549__A2 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net84 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net93 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3518__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3721__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3253__I mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ _1043_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5474__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5226__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ _2707_ _2733_ _2711_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4922_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _1862_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5908__I _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3804_ _0803_ _0828_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4784_ _1803_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _0156_ net115 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3735_ _0677_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3428__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6454_ mod.des.des_dout\[22\] net7 _3071_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3666_ _3215_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5162__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6385_ mod.des.des_dout\[11\] net9 _3027_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6632__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3597_ mod.registers.r14\[2\] _0624_ _0464_ mod.registers.r6\[2\] _0625_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5336_ _2237_ _2292_ _2297_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3712__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _2157_ _2251_ _2254_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4218_ _0908_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3476__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ mod.pc_2\[10\] _2178_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4149_ mod.funct3\[2\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6414__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4976__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6017__I1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4722__I _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4900__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3703__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3467__A1 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3467__B2 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6405__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6505__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6333__B _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6655__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3520_ _0419_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3451_ mod.registers.r2\[6\] _0477_ _0478_ mod.registers.r3\[6\] _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6170_ mod.des.des_dout\[20\] _2838_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3382_ mod.registers.r1\[7\] _3231_ _3234_ mod.registers.r13\[7\] _0410_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4300__C _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5121_ _2103_ _2127_ _2128_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _2037_ _2060_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _1028_ _1029_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_38_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _2714_ _2717_ _2718_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _1927_ _1928_ _1892_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5885_ mod.valid1 _2653_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4836_ _0730_ _0503_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4430__I0 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _1793_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5922__A3 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6506_ _0139_ net118 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3933__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3718_ _0739_ _0740_ _0741_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4698_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6437_ _3063_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5373__I _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3649_ _0435_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5686__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6368_ _3021_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3697__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3697__B2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ mod.registers.r3\[8\] _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _2086_ _2897_ _2972_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6486__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__A2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6528__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3621__B2 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5548__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6678__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5992__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3924__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5677__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3688__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3531__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout164_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _2491_ _2522_ _2527_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _1237_ _1646_ _1648_ _1193_ _1229_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5365__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4552_ _1412_ _1575_ _1576_ _1456_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3915__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3503_ mod.registers.r9\[5\] _0425_ _0429_ mod.registers.r10\[5\] _0531_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4483_ _0683_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3391__A3 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6222_ _0711_ _2924_ _2920_ mod.instr\[13\] _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3434_ mod.registers.r11\[6\] _3164_ _3167_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6153_ mod.des.des_dout\[15\] _2872_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3365_ _3215_ _3217_ _3209_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ mod.pc_1\[13\] _2820_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4479__I0 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3296_ mod.instr_2\[11\] mod.instr_2\[10\] _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _2039_ _2041_ _2050_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3441__I _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__S0 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__B1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4643__A3 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3851__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4981__B _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3851__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6820__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ mod.pc\[0\] _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3603__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__I0 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _2652_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4819_ _1739_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4159__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5799_ mod.registers.r13\[7\] _2605_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6199__I _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3685__A4 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_216 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_227 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_238 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6084__A2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_249 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3842__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5347__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5898__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6058__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4357__I _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6843__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6840_ _0067_ net183 mod.ldr_hzd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _0401_ net168 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4389__A2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3983_ _1007_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4092__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5722_ mod.registers.r11\[11\] _2556_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__B1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ mod.registers.r10\[0\] _2517_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5916__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _1352_ _1351_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5584_ _2379_ _2464_ _2467_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4010__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4010__B2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4535_ _1559_ _1560_ _1562_ _1181_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4561__A2 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3436__I _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _1147_ _1148_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4976__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6205_ _1710_ _2910_ _2913_ mod.instr\[7\] _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3417_ _0438_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5510__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _0874_ _1223_ _1423_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3521__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6136_ _2663_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3348_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A2 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ _2794_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3279_ _3131_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5018_ _0895_ _0900_ _1853_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5329__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4001__A1 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4001__B2 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3346__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4304__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4177__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4068__B2 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__A1 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__B2 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__B1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4240__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout127_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3256__I _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _1300_ _1308_ _1310_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_99_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4251_ _1271_ _1277_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5471__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3503__B1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4182_ _1208_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4059__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__I _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _0050_ net184 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _0384_ net186 mod.pc_1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3966_ mod.registers.r9\[13\] _0855_ _0863_ mod.registers.r1\[13\] _0994_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6739__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5705_ _2543_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6685_ _0318_ net102 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3897_ mod.registers.r5\[10\] _0487_ _0484_ mod.registers.r4\[10\] _0475_ mod.registers.r12\[10\]
+ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__3990__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _2474_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5731__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ mod.registers.r8\[7\] _2453_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4518_ _1360_ _1477_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _2382_ _2408_ _2412_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6287__A2 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _1037_ _0726_ _1231_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6119_ mod.instr\[7\] _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5798__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4725__I mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__C1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4222__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__D _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4773__A2 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6278__A2 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3264__A2 _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6202__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ mod.registers.r11\[9\] _0799_ _0786_ mod.registers.r5\[9\] _0848_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4213__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3751_ mod.pc_2\[8\] _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_9_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _3082_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3682_ _3179_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5421_ _2357_ _2347_ _2358_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5713__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _2138_ _2303_ _2309_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4303_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ _2245_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ _1258_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4165_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4096_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3589__C _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__S _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _0033_ net162 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4204__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ _3100_ _2013_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5952__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6737_ _0367_ net151 mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3949_ _0639_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4755__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3802__I1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6668_ _0301_ net135 mod.registers.r12\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ _2491_ _2484_ _2492_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4507__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _0232_ net74 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__B _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A2 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4746__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout70 net73 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout81 net84 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4190__I _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout92 net96 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3954__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3534__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout194_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _2730_ _2732_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1942_ _1943_ mod.pc\[5\] _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4985__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ _0608_ _0618_ _1849_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6187__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3803_ _0456_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4783_ _1758_ _1796_ _1799_ _1761_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3945__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6522_ _0155_ net117 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3734_ _0734_ _0735_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6453_ _3072_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3665_ _3202_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ _2144_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _3030_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3596_ _3183_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5335_ mod.registers.r3\[15\] _2293_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ mod.registers.r2\[5\] _2252_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4217_ _1238_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5197_ _2148_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3476__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4148_ _1175_ _3122_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4079_ _1082_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4425__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3936__B1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__I _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6350__A1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3467__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout207_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3450_ _3223_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6341__A1 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6341__B2 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3381_ _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ mod.registers.r1\[1\] _2118_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ _0957_ mod.funct7\[2\] _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4655__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4002_ mod.registers.r12\[12\] _0555_ _0865_ mod.registers.r2\[12\] _0859_ mod.registers.r3\[12\]
+ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_38_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__C1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ mod.pc\[1\] _2714_ _2711_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1833_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5884_ _2656_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _1860_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3439__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4766_ _0523_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4430__I1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3394__A1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6505_ _0138_ net119 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3717_ mod.registers.r13\[0\] _3233_ _3212_ mod.registers.r14\[0\] _0744_ _0745_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4697_ _3117_ _1723_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6436_ mod.des.des_dout\[14\] net17 _3061_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3648_ mod.pc_2\[3\] _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_106_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6367_ mod.des.des_dout\[3\] net19 _3017_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3579_ mod.registers.r1\[2\] _0483_ _0484_ mod.registers.r4\[2\] _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3697__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5318_ _2274_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6298_ mod.rd_3\[3\] _2962_ _2967_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5249_ _2090_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4249__I1 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3621__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3688__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4637__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5739__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5062__A1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout157_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3612__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3259__I _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4620_ _1246_ _1239_ _1647_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1278_ _1461_ _1544_ _1361_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3502_ mod.registers.r15\[5\] _0474_ _0475_ mod.registers.r12\[5\] _0530_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4482_ _1278_ _1509_ _1228_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5117__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6221_ _2796_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3433_ mod.registers.r5\[6\] _0460_ _3160_ mod.registers.r10\[6\] _0461_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6152_ _2663_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5103_ _2110_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _2814_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _3137_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4628__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4479__I1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ mod.pc_2\[11\] _2040_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__S1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3300__B2 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4643__A4 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3851__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6254__B _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _2701_ _2702_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3603__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4818_ mod.pc0\[0\] _1835_ _1841_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5356__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5798_ _2353_ _2604_ _2608_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4749_ _3221_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5384__I _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _2367_ _3048_ _3052_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput36 net36 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4867__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_217 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_228 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_239 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5559__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A2 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A1 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3542__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4086__A2 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__I _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6770_ _0400_ net173 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4389__A3 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3982_ _1009_ _1002_ _1005_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5721_ _2499_ _2555_ _2559_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3597__B2 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5338__A2 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4603_ _1427_ _1452_ _1485_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5583_ mod.registers.r8\[13\] _2465_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4534_ _1407_ _1410_ _1561_ _1511_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6518__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4465_ _0544_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3416_ _0440_ _0441_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6204_ _2903_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4396_ _0876_ _1217_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5510__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3521__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6135_ mod.instr\[11\] _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3521__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3347_ mod.instr_2\[17\] _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6668__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3452__I _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _2753_ _2803_ _2810_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3278_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5274__A1 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _2021_ _1348_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_45_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4283__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3588__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3588__B2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5919_ _2690_ _2691_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4785__B1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4001__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4068__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4407__B _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__A1 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6810__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4250_ _0621_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3503__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3503__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4181_ _1190_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4059__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6822_ _0049_ net182 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6753_ _0383_ net151 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3965_ mod.registers.r10\[13\] _0991_ _0992_ mod.registers.r13\[13\] _0993_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__I _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _2541_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6684_ _0317_ net134 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3896_ mod.registers.r15\[10\] _0474_ _0493_ mod.registers.r10\[10\] _0494_ mod.registers.r7\[10\]
+ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_109_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3990__A1 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3990__B2 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5635_ _2472_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3447__I _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5731__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5566_ _2354_ _2452_ _2456_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3742__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4479__S _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4517_ _1259_ _1260_ _1136_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__I _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5497_ mod.registers.r6\[14\] _2409_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6490__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4448_ _1473_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5495__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4379_ _1235_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6118_ _2847_ _2839_ _2849_ _2843_ _2844_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ mod.pc_1\[1\] _2797_ _2799_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__B1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4758__C2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3430__B1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5789__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__B _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4213__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ _0686_ _0773_ _0774_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ mod.registers.r6\[1\] _0572_ _0516_ mod.registers.r12\[1\] _0709_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3267__I mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ mod.registers.r5\[7\] _2348_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ mod.registers.r4\[3\] _2305_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5482__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4302_ _1329_ _1216_ _1284_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5282_ _2243_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4233_ _1259_ _1260_ _0726_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _3117_ _1117_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout52_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3660__B1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6805_ _0032_ net181 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ mod.pc0\[9\] _1887_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4204__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6856__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0366_ net153 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3948_ mod.registers.r4\[13\] _0974_ _0975_ mod.registers.r11\[13\] _0976_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5952__A2 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6667_ _0300_ net131 mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _0878_ _0763_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5618_ mod.registers.r9\[7\] _2485_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6598_ _0231_ net74 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5549_ _2443_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5392__I _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__I _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5468__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4515__I0 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4979__B1 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5995__C _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout71 net73 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout82 net84 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3954__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout93 net96 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__B2 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__CLK net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3550__I _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout187_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3890__B1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4434__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4920_ _1838_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6879__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _1653_ _1591_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_21_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4198__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3802_ _0658_ _0710_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4782_ _1800_ _1805_ _1808_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _0154_ net118 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3733_ _0747_ _0748_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3945__B2 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6452_ mod.des.des_dout\[21\] net6 _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3664_ mod.registers.r10\[1\] _0429_ _0548_ mod.registers.r11\[1\] _0692_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_134_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2343_ _2332_ _2344_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6383_ mod.des.des_dout\[10\] net8 _3027_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3595_ mod.registers.r8\[2\] _0457_ _3160_ mod.registers.r10\[2\] _0623_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4370__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5334_ _2231_ _2292_ _2296_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6111__A2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__I _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ _2145_ _2251_ _2253_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4216_ _1188_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5196_ _2176_ _2194_ _2195_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4673__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4147_ mod.funct3\[1\] _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3460__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4078_ _0413_ _1034_ _1035_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4425__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5387__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4291__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3936__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _0349_ net147 mod.pc0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3936__B2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3400__A3 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4361__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4113__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5861__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5613__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3475__I0 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3927__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout102_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _3232_ _3229_ _3207_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6551__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5050_ _2063_ _2051_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4655__A2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5852__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ mod.registers.r15\[12\] _0558_ _0898_ mod.registers.r6\[12\] _1029_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3458__A3 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__B1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__C2 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5604__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _2708_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__A2 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ mod.pc\[4\] _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5883_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _3111_ _3115_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ mod.instr_2\[4\] _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4979__C _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4430__I2 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _0137_ net72 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4591__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3716_ _0742_ _3208_ _0613_ _0614_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__3394__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _3112_ _3114_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6435_ _3062_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3455__I _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3647_ _0648_ _0656_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6332__A2 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _3020_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3578_ mod.registers.r7\[2\] _0494_ _0478_ mod.registers.r3\[2\] _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _2272_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6297_ _2970_ _2897_ _2971_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6096__A1 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _2099_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4286__I _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3854__B1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5179_ _2177_ _1986_ _2149_ _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6399__A2 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6006__I _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5845__I _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4582__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__C1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4334__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3688__A3 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__I _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4022__B1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4550_ _1236_ _1577_ _1454_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ mod.registers.r8\[5\] _0416_ _0420_ mod.registers.r11\[5\] _0529_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _1507_ _1508_ _1234_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4325__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6220_ _2651_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3432_ _3156_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6151_ mod.instr\[15\] _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3363_ mod.instr_2\[16\] _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5102_ _1860_ _3124_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _2055_ _2819_ _2821_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3294_ _3146_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5033_ _0000_ _1032_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3836__B1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3300__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ mod.pc0\[13\] _2678_ _2671_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _2650_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6270__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ mod.registers.r13\[6\] _2605_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4564__A1 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _1765_ _1775_ _0693_ _0413_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_5_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4679_ _1288_ _1348_ _1671_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_107_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ mod.registers.r15\[10\] _3049_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4867__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6349_ _3007_ _3009_ _2993_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5816__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_218 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_229 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A2 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__I _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5807__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3818__B1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6355__B _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3833__A3 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3981_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ mod.registers.r11\[10\] _2556_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3597__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ _2513_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4602_ _1517_ _1537_ _1574_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__4546__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _2374_ _2464_ _2466_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _1358_ _1409_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6299__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _1147_ _1148_ _1490_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6203_ _2907_ _2912_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3415_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4395_ _1303_ _1314_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6134_ _2859_ _2851_ _2861_ _2855_ _2856_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout82_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3521__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ mod.pc_1\[7\] _2805_ _2807_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3277_ _3121_ _3123_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3809__B1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ _3101_ _2031_ _2032_ _1997_ _2033_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_39_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6265__B _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5918_ _2683_ mod.pc0\[7\] _2684_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4785__A1 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4785__B2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ _2364_ _2637_ _2640_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6159__C _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__A2 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6762__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3579__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4423__B _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3553__I _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3503__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4317__C _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6205__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6205__B2 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6821_ _0048_ net180 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _0382_ net186 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4767__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3964_ _0480_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ _2481_ _2542_ _2548_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6683_ _0316_ net126 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3895_ mod.registers.r8\[10\] _0858_ _0859_ mod.registers.r3\[10\] _0923_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4519__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__B2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _2216_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3990__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5565_ mod.registers.r8\[6\] _2453_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6635__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4516_ _0684_ _0643_ _1368_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ _2379_ _2408_ _2411_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4447_ _1460_ _1245_ _1474_ _1371_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3463__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _1405_ _1295_ _1393_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6117_ mod.des.des_dout\[6\] _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ mod.registers.r4\[7\] _3177_ _3181_ mod.registers.r2\[7\] _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6048_ _2710_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4294__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__B2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__A3 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3430__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3430__B2 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3733__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3373__I _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A2 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3249__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6508__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3421__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__I _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout132_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3680_ mod.registers.r8\[1\] _0581_ _0576_ mod.registers.r13\[1\] _0708_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5174__A1 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _2133_ _2303_ _2308_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3724__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _1215_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5281_ _2209_ _2257_ _2262_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5477__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _1132_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ _1188_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6426__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _1114_ _1115_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5003__I _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout45_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3660__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__B2 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6804_ _0031_ net181 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4996_ _2014_ _1928_ _1892_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _0365_ net152 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3947_ _0626_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _0299_ net133 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3878_ _0890_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5165__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _2173_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6597_ _0230_ net46 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4912__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5479_ mod.registers.r6\[7\] _2397_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5468__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4515__I1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4140__A2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6417__A1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4979__B2 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6800__CLK net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6172__C _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net68 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout72 net73 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3954__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3706__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3831__I _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3890__A1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3890__B2 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3987__B _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3642__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__I _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3642__B2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3801_ _0445_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4198__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3278__I _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ mod.instr_2\[6\] _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6520_ _0153_ net69 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3945__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3732_ mod.pc_2\[0\] _0507_ _0753_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _3060_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3663_ mod.registers.r8\[1\] _0416_ _0425_ mod.registers.r9\[1\] _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_109_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5402_ mod.registers.r5\[3\] _2334_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5698__A2 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6382_ _3029_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3594_ mod.pc_2\[2\] _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5333_ mod.registers.r3\[14\] _2293_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4370__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ mod.registers.r2\[4\] _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4215_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5195_ mod.registers.r1\[9\] _2185_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4146_ _1125_ _1172_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3881__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4077_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4433__I0 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _3101_ _1995_ _1996_ _1997_ _1998_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6718_ _0348_ net148 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3936__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _0282_ net123 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4521__B _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A2 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4113__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4664__A3 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__I1 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3927__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6358__B _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4000_ mod.registers.r5\[12\] _0819_ _0858_ mod.registers.r8\[12\] _1028_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3863__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__B2 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _1869_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4606__B _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _3105_ _1726_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_80_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ _2662_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5368__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _1072_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4764_ _1784_ _1787_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6503_ _0136_ net72 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3715_ mod.registers.r15\[0\] _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4430__I3 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _3119_ _1711_ _1715_ _1719_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6434_ mod.des.des_dout\[13\] net16 _3061_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3646_ _0455_ _0660_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6365_ mod.des.des_dout\[2\] net18 _3017_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5540__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3577_ _0451_ _0505_ _0595_ _0603_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_114_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _2174_ _2280_ _2285_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ mod.rd_3\[2\] _2962_ _2967_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6268__B _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__A2 _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _2239_ _2096_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3471__I _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _0833_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3854__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3854__B2 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _0600_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6719__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6022__I mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3790__C2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3381__I _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__A1 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4270__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4022__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4022__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5770__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout212_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3500_ mod.registers.r13\[5\] _3234_ _3213_ mod.registers.r14\[5\] _0528_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3781__B1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4480_ _1155_ _1249_ _1265_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4325__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3431_ mod.registers.r13\[6\] _3140_ _3144_ mod.registers.r1\[6\] _0459_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5522__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ _2871_ _2863_ _2873_ _2867_ _2868_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3362_ _3200_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ mod.ins_ldr_3 mod.valid_out3 net15 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ mod.pc_1\[12\] _2820_ _2815_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3291__I _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3293_ mod.instr_2\[13\] _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3836__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__B2 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _2689_ _2068_ _2071_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_34_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ _2649_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6002__A2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4816_ _1843_ _1833_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _2350_ _2604_ _2607_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5210__B1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4564__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _0427_ _0695_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3466__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _1691_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6417_ _2364_ _3048_ _3051_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4498__S _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _3215_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5513__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5681__I _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput27 net27 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput38 net38 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__B1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6348_ _2997_ _1812_ _3008_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4297__I _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ mod.valid_out3 _2091_ _2657_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_219 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5752__A1 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6691__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3818__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout162_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ mod.pc_2\[13\] _3127_ _0970_ _0983_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4794__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ _1591_ _1607_ _1611_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__A1 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5581_ mod.registers.r8\[12\] _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4546__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4532_ _1416_ _1541_ _1456_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6299__A2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _0451_ _0505_ _0604_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3506__B1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6202_ _1809_ _2910_ _2904_ mod.instr\[6\] _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3414_ mod.funct3\[2\] _0437_ _3124_ mod.instr_2\[1\] _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4394_ _1186_ _1419_ _1421_ _1330_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6133_ mod.des.des_dout\[10\] _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3345_ _3197_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout75_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _2746_ _2803_ _2809_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3276_ _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3809__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3809__B2 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5015_ _3092_ _2022_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4482__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6564__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4234__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _2689_ _1977_ _1980_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5982__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3588__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5848_ mod.registers.r14\[9\] _2638_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4537__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4225__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6210__I _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6150__B2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6205__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _0047_ net182 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _0493_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6751_ _0381_ net186 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4767__A2 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ mod.registers.r11\[3\] _2544_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6682_ _0315_ net133 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3894_ _0911_ _0569_ _0916_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4519__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _2501_ _2494_ _2502_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5564_ _2351_ _2452_ _2455_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4515_ _0597_ _0473_ _0593_ _1439_ _1265_ _1204_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5495_ mod.registers.r6\[13\] _2409_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3742__A3 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__I _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _1149_ _1259_ _1260_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6116_ _2825_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3328_ _3180_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6047_ _2703_ _2795_ _2798_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3259_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4455__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__B1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3430__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__A1 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__A3 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3249__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3709__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4300_ _1325_ _1253_ _1327_ _1186_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_5_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5280_ mod.registers.r2\[11\] _2258_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _1131_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4093_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4437__A1 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4988__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ _0030_ net180 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ mod.pc\[9\] _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__I mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3948__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6602__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6734_ _0364_ net153 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3946_ _0628_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3877_ _0901_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6665_ _0298_ net132 mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5616_ _2489_ _2484_ _2490_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5165__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _0229_ net56 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4912__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5547_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5478_ _2354_ _2396_ _2400_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4429_ _1453_ _1455_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4515__I2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6417__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4428__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3649__I _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout40 net50 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net55 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4061__C1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout62 net67 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout73 net78 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6353__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A3 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4667__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3890__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6625__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ _0804_ _0815_ _0826_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4780_ mod.instr_2\[5\] _1806_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5395__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3731_ _0754_ _0755_ _0757_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6450_ _3070_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3662_ mod.registers.r6\[1\] _0418_ _3223_ mod.registers.r3\[1\] _0430_ mod.registers.r7\[1\]
+ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6381_ mod.des.des_dout\[9\] net7 _3027_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3593_ _0619_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5332_ _2225_ _2292_ _2295_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _2245_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4214_ _0621_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5194_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3330__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4145_ _1112_ _1076_ _1171_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_29_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _0539_ _1103_ _3196_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__I _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4978_ _1873_ _1517_ _3098_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4433__I1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6717_ _0347_ net184 mod.valid1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3929_ mod.pc_2\[13\] _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _0281_ net80 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5138__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _0212_ net52 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4897__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4649__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3932__I _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5310__A2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6648__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3927__A3 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5129__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout192_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3863__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5769__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5065__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5950_ _1855_ _1829_ _1866_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_52_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4901_ _1728_ _1923_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ mod.valid0 _2653_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4832_ _1858_ _1573_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__B1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4763_ _1789_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _0135_ net69 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3714_ mod.registers.r12\[0\] _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6317__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4694_ _1710_ _1721_ _1312_ _1713_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4341__C _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3645_ mod.pc_2\[3\] _0661_ _0666_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6364_ _3019_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3576_ _3193_ _0450_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3551__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ mod.registers.r3\[7\] _2281_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3752__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6295_ _0440_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ _2091_ _2094_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5177_ _2106_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3854__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _1155_ _0450_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__A1 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input18_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ mod.registers.r9\[15\] _0977_ _0968_ mod.registers.r10\[15\] _1087_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5359__A2 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6308__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3790__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B2 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__A2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__I _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__I _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4022__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5770__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3781__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3781__B2 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6813__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3430_ mod.registers.r8\[6\] _0457_ _3152_ mod.registers.r9\[6\] _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout205_I net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3361_ mod.registers.r15\[7\] _3206_ _3210_ mod.registers.r12\[7\] _3213_ mod.registers.r14\[7\]
+ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_98_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ _2108_ _1733_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _2804_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3292_ mod.registers.r13\[7\] _3140_ _3144_ mod.registers.r1\[7\] _3145_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5286__A1 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A2 _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _2021_ _1652_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3836__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _2699_ _2700_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ net11 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5210__A1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ mod.registers.r13\[5\] _2605_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6123__I mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4746_ _1399_ _1072_ _1740_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4564__A3 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5761__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4677_ _1402_ _1695_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6493__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ mod.registers.r15\[9\] _3049_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3628_ _0649_ _0650_ _0651_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5513__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A1 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3524__B2 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6347_ _2086_ _2965_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3559_ mod.registers.r7\[4\] _0585_ _0586_ mod.registers.r12\[4\] _0587_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _2092_ _2896_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5277__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5229_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6836__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3515__A1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3392__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5268__A1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3818__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__B1 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout155_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3451__B1 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4794__A3 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4600_ _1504_ _1619_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5580_ _2446_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _1555_ _1558_ _1228_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5782__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4462_ _1145_ _1443_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3506__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ _2907_ _2911_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3413_ _3217_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4393_ _1377_ _1378_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6132_ _2825_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3344_ _3110_ _3113_ mod.instr_2\[1\] _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ _3116_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6063_ mod.pc_1\[6\] _2805_ _2807_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3809__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5014_ _0926_ _0930_ _1853_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6709__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout68_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4482__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5431__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _2677_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6859__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3442__B1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _2359_ _2637_ _2639_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3993__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5778_ _2100_ _2567_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _1753_ _1754_ _1755_ _1756_ _1749_ _1750_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_135_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5498__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__I _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5670__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3681__B1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__I _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4704__C _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3984__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5088__B _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5489__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6150__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5107__I _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3850__I mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A2 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5413__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _0380_ net187 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ mod.registers.r12\[13\] _0893_ _0823_ mod.registers.r2\[13\] _0990_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5964__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5701_ _2479_ _2542_ _2547_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6681_ _0314_ net133 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3893_ _0917_ _0918_ _0919_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5632_ mod.registers.r9\[11\] _2495_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5716__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3727__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5563_ mod.registers.r8\[5\] _2453_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4514_ _1119_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5494_ _2374_ _2408_ _2410_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4445_ _1273_ _1245_ _1472_ _1244_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6531__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4376_ _1399_ _1215_ _3129_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_59_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6115_ mod.instr\[6\] _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3327_ _3178_ _3179_ _3142_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ mod.pc_1\[0\] _2797_ _2751_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3258_ _3110_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__A2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6681__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3663__B1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__C _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3966__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3966__B2 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _0106_ net202 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__I _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4391__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4766__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5597__I _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A2 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3957__A1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3709__A1 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6221__I _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ _1003_ _1196_ _1136_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _0780_ _0765_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3645__B1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_370 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _0029_ net170 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4994_ _2001_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3948__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ _0363_ net149 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ mod.registers.r8\[13\] _0971_ _0972_ mod.registers.r2\[13\] _0973_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _0297_ net79 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3876_ _0545_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5615_ mod.registers.r9\[6\] _2485_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6595_ _0228_ net89 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6131__I mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5546_ _2300_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3581__C1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6114__A2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ mod.registers.r6\[6\] _2397_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4125__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4428_ _0775_ _1184_ _1123_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4515__I3 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4359_ _1162_ _1169_ _1351_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3490__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__B1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _2756_ _2774_ _2779_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_73_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__B1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4535__B _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4254__C _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6050__A1 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4061__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout41 net42 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4600__A2 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net55 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout63 net64 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout74 net77 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout96 net97 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4270__B _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6041__I _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4364__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A2 _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__I _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5616__A1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__B1 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4445__B _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ mod.registers.r9\[0\] _0639_ _0582_ mod.registers.r3\[0\] _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3661_ _0687_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4355__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5400_ _2137_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6380_ _3028_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3592_ _3108_ _0444_ _0500_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_115_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ mod.registers.r3\[13\] _2293_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ _2243_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4658__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _1239_ _1046_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ mod.des.des_dout\[30\] _2187_ _2189_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_69_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3866__B1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ _1076_ _1171_ _1112_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3881__A3 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4075_ mod.registers.r12\[15\] _0893_ _1098_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_55_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3618__B1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout50_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6126__I _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _3094_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5965__I mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__I2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6716_ _0346_ net189 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3928_ _0946_ _0953_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6647_ _0280_ net79 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ mod.registers.r5\[11\] _0786_ _0792_ mod.registers.r2\[11\] _0887_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6578_ _0211_ net51 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4897__A2 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _2365_ _2429_ _2432_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4649__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5846__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3434__B _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__B1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__B1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4337__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4888__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3545__C1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5837__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3344__B mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6262__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6742__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4900_ _1736_ _1914_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ _2093_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6014__A1 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _1309_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4025__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6892__CLK net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__B2 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1756_ _1777_ _1778_ _1753_ _1779_ _1755_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_119_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _0134_ net70 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ mod.registers.r8\[0\] _0415_ _0419_ mod.registers.r11\[0\] _0741_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4693_ _1113_ _1720_ _1717_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6317__A2 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4328__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6432_ mod.des.des_counter\[2\] _2074_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ _0667_ _0668_ _0669_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ mod.des.des_dout\[1\] net17 _3017_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3575_ _0598_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ _2167_ _2280_ _2284_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3551__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _1797_ _2897_ _2969_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5828__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _2211_ _2237_ _2238_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3303__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ _2106_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4864__I _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4127_ _0597_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5056__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ mod.registers.r6\[15\] _0960_ _0978_ mod.registers.r12\[15\] _1086_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6005__A1 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5695__I _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6308__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4104__I _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3790__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3943__I _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5819__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__CLK net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__A1 _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4949__I _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _3212_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _1966_ _2034_ _2035_ _1997_ _2046_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3297__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5038__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6235__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ _2670_ mod.pc0\[12\] _2671_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5863_ _2384_ _2643_ _2648_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4549__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _1836_ _1838_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5794_ _2345_ _2604_ _2606_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _1752_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6638__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4676_ _1309_ _1296_ _1692_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6010__I1 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6415_ _2359_ _3048_ _3050_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3627_ mod.registers.r13\[3\] _3234_ _3213_ mod.registers.r14\[3\] _0654_ _0655_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3763__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput29 net29 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3524__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6346_ _1745_ _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3558_ _3189_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _0957_ _2893_ _2958_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3489_ mod.registers.r7\[5\] _0467_ _0516_ mod.registers.r12\[5\] _0517_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_76_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ mod.des.des_dout\[34\] _2152_ _2221_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_97_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5159_ _3109_ _3165_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__C _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4960__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4769__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3515__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5268__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4009__I _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3451__A1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3451__B2 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A4 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout148_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4251__I0 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4530_ _1191_ _1556_ _1557_ _1236_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4461_ _1272_ _1150_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6200_ _2909_ _2910_ _2904_ mod.instr\[5\] _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3506__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ mod.instr_2\[5\] _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4392_ _1243_ _1370_ _1256_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6131_ mod.instr\[10\] _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _3195_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2742_ _2803_ _2808_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3274_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _2018_ _2020_ _2030_ _2001_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A1 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5915_ _2687_ _2688_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3758__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3442__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3442__B2 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ mod.registers.r14\[8\] _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3993__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__A1 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _2511_ _2589_ _2594_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4728_ mod.ldr_hzd\[3\] _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3707__B _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4659_ _1076_ _1320_ _1686_ _3131_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6329_ _2994_ _2995_ _2993_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4170__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__I _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3681__B2 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3433__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3433__B2 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3984__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__I _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3736__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ mod.registers.r7\[13\] _0987_ _0988_ mod.registers.r11\[13\] _0989_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4472__I0 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ mod.registers.r11\[2\] _2544_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ _0313_ net82 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3892_ mod.registers.r4\[10\] _0570_ _0799_ mod.registers.r11\[10\] _0920_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ _2208_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4924__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3727__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _2346_ _2452_ _2454_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4513_ _1453_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5493_ mod.registers.r6\[12\] _2409_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4202__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4444_ _1263_ _1259_ _1260_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _1125_ _1397_ _1398_ _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_98_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6429__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _2845_ _2839_ _2846_ _2843_ _2844_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout80_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ _3158_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3257_ mod.instr_2\[2\] _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6826__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3663__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3663__B2 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5189__B _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3488__I _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3966__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _0105_ net198 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5168__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _2336_ _2624_ _2628_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4391__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4112__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5878__I _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3709__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4134__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__A1 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6849__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_360 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3645__B2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_371 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4692__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6801_ _0028_ net171 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5398__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _1879_ _1999_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3948__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3944_ _0571_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6732_ _0362_ net152 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6663_ _0296_ net79 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3875_ _3147_ _0829_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6412__I _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5614_ _2166_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ _0227_ net58 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5545_ _2085_ _2441_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3581__B1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3581__C2 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5476_ _2351_ _2396_ _2399_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _1093_ _1200_ _1454_ _1361_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5322__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4125__A2 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3771__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__B1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4358_ _1126_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3884__B2 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3309_ _3133_ _3158_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4289_ _1311_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _2777_ _2763_ _2782_ _2741_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3636__B2 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3720__B _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4061__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout42 net49 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4061__B2 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout75 net77 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3946__I _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout86 net140 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net101 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3627__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__B2 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5401__I _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4445__C _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6521__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout130_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__I _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3660_ mod.registers.r5\[1\] _0487_ _0477_ mod.registers.r2\[1\] _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4355__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3591_ _0546_ _0608_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6671__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5330_ _2217_ _2292_ _2294_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5261_ _2138_ _2244_ _2250_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5304__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4212_ _1131_ _1132_ _1008_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4658__A3 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _2113_ _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3866__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3866__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4143_ _1128_ _1170_ _1078_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3330__A3 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4074_ _1099_ _1100_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__B _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3618__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__C _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout43_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__A2 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4043__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ _0815_ _0826_ _1915_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4433__I3 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6715_ _0002_ _0006_ net201 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3927_ _0954_ _0901_ _0904_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3766__I _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6142__I _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3858_ mod.registers.r4\[11\] _0570_ _0799_ mod.registers.r11\[11\] _0886_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6646_ _0279_ net80 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5543__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6577_ _0210_ net52 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5981__I mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3789_ _3234_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ mod.registers.r7\[9\] _2430_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6298__B _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5459_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4729__S0 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net213 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3857__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__B2 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3609__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3609__B2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__I _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6544__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A2 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__B2 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6694__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5891__I _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3545__B1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3545__C2 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__C1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3848__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A3 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout178_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4025__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__B2 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4576__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _1754_ _1775_ _1788_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6500_ _0133_ net43 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3784__B1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3712_ mod.registers.r9\[0\] _0424_ _0428_ mod.registers.r10\[0\] _0740_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _1288_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4328__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6431_ _2384_ _3054_ _3059_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3643_ mod.registers.r13\[3\] _3139_ _3143_ mod.registers.r1\[3\] _0670_ _0671_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6362_ _3018_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _0600_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ mod.registers.r3\[6\] _2281_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6293_ mod.rd_3\[1\] _2962_ _2967_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4210__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5244_ mod.registers.r1\[15\] _2218_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5175_ _2102_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _1129_ _1144_ _1146_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_110_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4366__B _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _1083_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ mod.pc0\[7\] _1909_ _1961_ _1979_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3775__B1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5516__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _0262_ net83 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4276__B _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6244__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4558__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__I _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3290_ _3134_ _3136_ _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _2689_ _2054_ _2057_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_19_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ mod.registers.r14\[15\] _2644_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5793_ mod.registers.r13\[4\] _2605_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3757__B1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _0712_ _1757_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4675_ _1334_ _1697_ _1699_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6414_ mod.registers.r15\[8\] _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3626_ _0652_ _3208_ _0613_ _0614_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3557_ _0467_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6345_ _2973_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6276_ mod.pc_1\[13\] _2665_ _2955_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _3189_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5227_ _2113_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4485__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5158_ _0452_ _2129_ _2148_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ _1131_ _1132_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_45_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ mod.rd_3\[0\] _2083_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5985__A1 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4960__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3903__B _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6882__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3451__A2 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4251__I1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4951__A2 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout210_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _0605_ _0778_ _1160_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3411_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4391_ _1262_ _1192_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6130_ _2857_ _2851_ _2858_ _2855_ _2856_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3342_ _3194_ _3124_ _3107_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ mod.pc_1\[5\] _2805_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3273_ _3125_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5012_ _1985_ _2022_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4219__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5914_ _2683_ mod.pc0\[6\] _2684_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6605__CLK net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3442__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ _2625_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ mod.registers.r12\[15\] _2590_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6755__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4727_ mod.ldr_hzd\[2\] _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4658_ _1059_ _1071_ _1073_ _1218_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _0612_ _0634_ _3188_ _0636_ _0615_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4589_ _1205_ _1616_ _1541_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6328_ _2909_ _2983_ _2978_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _2657_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3949__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6325__I _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3433__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4481__I1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5186__A2 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4449__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__S _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6628__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A2 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _0548_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__I1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6778__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3891_ mod.registers.r8\[10\] _0791_ _0797_ mod.registers.r10\[10\] _0919_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ _2499_ _2494_ _2500_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ mod.registers.r8\[4\] _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ _1511_ _1502_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5492_ _2390_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _1468_ _1157_ _0601_ _1180_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4374_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3896__C1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ mod.des.des_dout\[5\] _2835_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3325_ _3157_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3256_ _3108_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6044_ _2793_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3663__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3769__I _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4612__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ _0104_ net206 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5828_ mod.registers.r14\[1\] _2626_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5759_ _2571_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4915__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6117__A1 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4549__B _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3654__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6055__I _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A1 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3406__A2 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__I _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__A1 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6004__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__I _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__B _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3342__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _3117_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_350 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__A1 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3645__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_361 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_372 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6800_ _0027_ net169 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _2004_ _2009_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6731_ _0361_ net141 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3943_ _0581_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6662_ _0295_ net80 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6347__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3874_ mod.funct7\[2\] _0869_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _2487_ _2484_ _2488_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _0226_ net57 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5544_ _2089_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3581__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5475_ mod.registers.r6\[5\] _2397_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _1183_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6370__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4369__B _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__I0 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__B1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__B2 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4357_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3884__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3308_ mod.registers.r5\[7\] _3156_ _3160_ mod.registers.r10\[7\] _3161_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4288_ _0954_ _0905_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5979__I _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3239_ net141 _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6027_ _2780_ _2781_ _2739_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__A2 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4061__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout43 net49 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net55 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout76 net77 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout87 net90 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_6_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5313__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6361__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3627__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4037__C1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6816__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ _0609_ _0610_ _0611_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5552__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5304__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ mod.registers.r2\[3\] _2246_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3315__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4211_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5191_ _1919_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3866__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4142_ _1162_ _1169_ _1011_ _1041_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ mod.registers.r2\[15\] _0823_ _0811_ mod.registers.r3\[15\] _1101_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3618__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _1984_ _1994_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5240__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _0001_ _0005_ net201 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__6423__I _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3926_ _0890_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6645_ _0278_ net81 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5039__I mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3857_ mod.registers.r7\[11\] _0585_ _0586_ mod.registers.r12\[11\] _0885_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6496__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6576_ _0209_ net91 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3788_ _0418_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _2360_ _2429_ _2431_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3782__I _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5458_ _2241_ _2299_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4729__S1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4409_ _1433_ _1435_ _1436_ _1430_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xfanout200 net215 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout211 net212 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5389_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3857__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5059__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3609__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4034__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6839__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3545__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3545__B2 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4742__C2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5470__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4025__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _0657_ _0693_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5773__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3784__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3711_ mod.registers.r5\[0\] _0422_ _3225_ mod.registers.r2\[0\] _0417_ mod.registers.r6\[0\]
+ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__3784__B2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4691_ _1710_ _1718_ _1712_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6430_ mod.registers.r15\[15\] _3055_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3642_ _0652_ _3175_ _3188_ _0636_ _0653_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6361_ mod.des.des_dout\[0\] net16 _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3573_ _0599_ _0498_ _0504_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5312_ _2157_ _2280_ _2283_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6292_ _1794_ _2819_ _2968_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5289__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5243_ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ _2140_ _2174_ _2175_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3551__B _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4125_ _1147_ _1148_ _1151_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ mod.registers.r7\[15\] _0962_ _0967_ mod.registers.r5\[15\] _1084_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3777__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5764__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3775__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3775__B2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3909_ _0931_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4889_ _1876_ _1897_ _1898_ _1852_ _1913_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6628_ _0261_ net66 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5516__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4575__I0 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6559_ _0192_ net92 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4557__B _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5407__I _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4311__I _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5691__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout190_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _2696_ _2698_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3454__B1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _2381_ _2643_ _2647_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4812_ _1837_ _1839_ mod.pc\[0\] _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5746__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5792_ _2598_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3757__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3757__B2 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ _1760_ _1764_ _1766_ _1770_ _0437_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4930__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4674_ _1230_ _1584_ _1701_ _1331_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3509__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6413_ _3036_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3625_ mod.registers.r15\[3\] _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5317__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4221__I _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4182__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _2999_ _3005_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3556_ mod.registers.r8\[4\] _0581_ _0582_ mod.registers.r3\[4\] _0583_ mod.registers.r5\[4\]
+ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6275_ _2062_ _2893_ _2957_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3487_ mod.registers.r4\[5\] _3177_ _3181_ mod.registers.r2\[5\] _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _1987_ _2110_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6148__I _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6684__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _2120_ _1951_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3693__B1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _1133_ _0932_ _1134_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5088_ _2091_ _2094_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input16_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4891__I _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4039_ mod.registers.r15\[14\] _0810_ _0811_ mod.registers.r3\[14\] _1067_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3987__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__I1 _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4306__I _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3739__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3410_ _0437_ _3197_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout203_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1344_ _1413_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3341_ mod.funct7\[2\] _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _2710_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ _3107_ _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A1 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ _1932_ _2025_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4925__B _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4219__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5967__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__I _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3978__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _2675_ _1960_ _1964_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6893_ _0120_ net200 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__I1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4216__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5844_ _2623_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5719__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ _2509_ _2589_ _2593_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4726_ mod.ldr_hzd\[1\] _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4657_ _1230_ _1465_ _1684_ _1301_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4155__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ _3174_ _0635_ _3134_ _3179_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4588_ _1266_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ _1768_ _2988_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3539_ _0545_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _0453_ _2940_ _2946_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4458__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5209_ _2104_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _2899_ _2902_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4449__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4472__I2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout153_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__S _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ mod.registers.r3\[10\] _0782_ _0586_ mod.registers.r12\[10\] _0918_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _2446_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4511_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5491_ _2388_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4442_ _1329_ _0600_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3896__B1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3896__C2 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6112_ mod.instr\[5\] _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3324_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5637__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3255_ _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4860__A2 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6062__A1 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6722__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__B1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _0103_ net206 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__B1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ _2328_ _2624_ _2627_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3785__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6872__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _2569_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _1734_ _1735_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5689_ mod.registers.r10\[15\] _2535_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4128__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3734__B _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4679__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5505__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4851__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3406__A3 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6071__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__A2 _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5415__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3342__A2 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5619__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6292__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6745__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__B _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_340 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_351 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_362 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4842__A2 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__B1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4991_ _2004_ _2009_ _1900_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _0360_ net141 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3942_ _0961_ _0964_ _0966_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _0294_ net81 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3873_ _0804_ _0895_ _0900_ _0827_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6347__A2 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5612_ mod.registers.r9\[5\] _2485_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6592_ _0225_ net93 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5543_ _2385_ _2435_ _2440_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5474_ _2346_ _2396_ _2398_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _1109_ _0775_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3869__B1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__A2 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__B2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__I1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _1182_ _1366_ _1375_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3307_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4287_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6026_ _2771_ _2775_ _2779_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3238_ _3092_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout44 net45 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout55 net62 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6859_ _0086_ net102 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout66 net67 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout77 net78 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout88 net90 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout99 net101 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6618__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5849__A1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__B1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__C2 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _1206_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5190_ _2110_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ _0909_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ mod.registers.r15\[15\] _0810_ _0898_ mod.registers.r6\[15\] _1100_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4028__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4974_ _1891_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6713_ _0000_ _0004_ net201 mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_3925_ _0947_ _0950_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _0277_ net63 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3856_ mod.registers.r9\[11\] _0781_ _0794_ mod.registers.r1\[11\] _0884_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6575_ _0208_ net92 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ _0807_ _0809_ _0812_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5526_ mod.registers.r7\[8\] _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4751__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5457_ _2385_ _2375_ _2386_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4503__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _0770_ _0771_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xfanout201 net215 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5388_ _2330_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout212 net213 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3711__C1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _1256_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5059__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ mod.pc\[9\] _2012_ _1842_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4562__C _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__A2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6192__B1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3545__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__B2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__A3 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3922__B _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6247__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4309__I _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5470__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4044__I _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6460__S _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3710_ _0736_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3784__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4981__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _1113_ _1708_ _3119_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3641_ mod.registers.r9\[3\] _3151_ _3170_ mod.registers.r3\[3\] _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3883__I mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4584__I1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3572_ _0498_ _0504_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ mod.registers.r3\[5\] _2281_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ mod.rd_3\[0\] _2820_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5242_ mod.des.des_dout\[36\] _2159_ _2233_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ mod.registers.r1\[7\] _2146_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5603__I _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4124_ _1149_ _1150_ _0776_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4055_ mod.registers.r1\[15\] _0965_ _0963_ mod.registers.r3\[15\] _1083_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5213__A2 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4957_ _1942_ _1943_ mod.pc\[7\] _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__S _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3908_ _0932_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4888_ _1899_ _1908_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3839_ _0862_ _0864_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6627_ _0260_ net67 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3793__I _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6558_ _0191_ net95 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _2337_ _2416_ _2420_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6489_ _0122_ net116 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4557__C _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4129__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__B _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6401__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A1 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6012__C _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4748__B _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5423__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__C _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout183_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3454__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3454__B2 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5860_ mod.registers.r14\[14\] _2644_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _2596_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3757__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _1767_ _3184_ _1762_ _1768_ _1769_ _0634_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4673_ _1325_ _1679_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6412_ _3034_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3624_ mod.registers.r12\[3\] _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3509__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _1761_ _3000_ _3001_ _2986_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4182__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3555_ _3156_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6274_ mod.pc_1\[12\] _2665_ _2955_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3486_ mod.registers.r3\[5\] _3171_ _0464_ mod.registers.r6\[5\] _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4658__B _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _2107_ _2060_ _2196_ _2220_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6829__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5156_ _2110_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3693__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__B2 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ _0754_ _0755_ _0757_ _0758_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _1797_ _2082_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4038_ mod.registers.r14\[14\] _0821_ _0988_ mod.registers.r11\[14\] _1066_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6482__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3788__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3996__A2 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5989_ _1960_ _1962_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3748__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__A1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__I _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3684__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4308__S0 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3698__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3987__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A1 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5418__I _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3340_ mod.pc_2\[7\] _3127_ _3192_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3271_ mod.instr_2\[2\] mod.instr_2\[0\] _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5153__I _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _2026_ _2027_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3675__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _2669_ _1947_ _2686_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3978__A2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3401__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _0119_ net203 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _2356_ _2631_ _2636_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ mod.registers.r12\[14\] _2590_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6501__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4725_ mod.ldr_hzd\[0\] _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5328__I _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4232__I _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4656_ _1683_ _1362_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3607_ _3137_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4155__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _1326_ _1612_ _1614_ _1511_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6326_ _2991_ _2992_ _2993_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3538_ _0546_ _0553_ _0561_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_115_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ mod.pc_1\[6\] _2941_ _2942_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3469_ _3195_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4458__A3 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _1953_ _2148_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6188_ _3111_ _2900_ _2891_ mod.instr\[2\] _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5998__I _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3666__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5139_ mod.des.des_dout\[25\] _2141_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_29_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3418__A1 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__B1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3311__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3981__I _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5646__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3657__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6524__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4472__I3 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout146_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5582__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__I _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4052__I _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4510_ _0761_ _1512_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5490_ _2371_ _2402_ _2407_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4441_ _1329_ _1468_ _1220_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5334__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4372_ _1399_ _1312_ _1178_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3896__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _2841_ _2839_ _2842_ _2843_ _2844_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3323_ _3174_ _3155_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5637__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3254_ _3106_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__B _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__I _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout59_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6062__A2 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4073__B2 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4612__A3 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ _0102_ net206 mod.des.des_dout\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3820__B2 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6442__I _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5826_ mod.registers.r14\[0\] _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _2491_ _2577_ _2582_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _1727_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5688_ _2509_ _2534_ _2538_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4128__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _1158_ _1319_ _1223_ _1156_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4679__A3 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3887__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _2659_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6547__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4137__I _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3811__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5013__B1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3925__B _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3878__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6020__C _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__B1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__A2 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_330 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_341 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_352 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_363 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4990_ _2007_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4055__B2 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ mod.registers.r5\[13\] _0967_ _0968_ mod.registers.r10\[13\] _0969_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ _0293_ net54 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3872_ _0896_ _0897_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5611_ _2156_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5555__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _0224_ net92 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5542_ mod.registers.r7\[15\] _2436_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5473_ mod.registers.r6\[4\] _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5606__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4424_ _1290_ _1446_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__B2 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ _1007_ _1223_ _1376_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4381__I2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3306_ _3146_ _3148_ _3157_ _3158_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6283__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _2771_ _2775_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3237_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4385__C _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3796__I _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout45 net48 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6858_ _0085_ net102 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout56 net57 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout67 net68 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout78 net85 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ mod.registers.r13\[11\] _2611_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5546__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout89 net97 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6789_ _0016_ net160 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6274__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4285__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__B2 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5537__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6458__S _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4140_ _1164_ _1167_ _0906_ _0938_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__B _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__A2 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ mod.registers.r5\[15\] _0819_ _0813_ mod.registers.r8\[15\] _1099_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4276__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4028__A1 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4028__B2 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5776__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _1985_ _1986_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6712_ _0345_ net74 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3924_ _0951_ _0937_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5528__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ _0276_ net87 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3855_ _0879_ _0880_ _0881_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3786_ mod.registers.r8\[8\] _0813_ _0551_ mod.registers.r7\[8\] _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6574_ _0207_ net91 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _2417_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4751__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5456_ mod.registers.r5\[15\] _2376_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4503__A2 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4407_ _1130_ _1434_ _1258_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5700__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout202 net203 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout213 net214 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3711__B1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4338_ _1344_ _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3711__C2 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__A2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4269_ _0946_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5071__I _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6008_ _2757_ _2760_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6192__A1 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__A2 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6885__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4981__A2 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ mod.registers.r7\[3\] _3187_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6183__A1 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ mod.pc_2\[6\] _3126_ _0463_ _0471_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5156__I _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3941__B1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _2145_ _2280_ _2282_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _2709_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _2190_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5172_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4123_ _1149_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4054_ _1003_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout41_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__I _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _1855_ _1829_ _1976_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6758__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3907_ _0869_ _0541_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ mod.pc0\[3\] _1909_ _1845_ _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_20_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6626_ _0259_ net66 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3838_ mod.registers.r2\[9\] _0865_ _0547_ mod.registers.r10\[9\] mod.registers.r14\[9\]
+ _0820_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5921__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _0190_ net88 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4724__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _3159_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5508_ mod.registers.r7\[1\] _2418_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6488_ _0121_ _0003_ net201 mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _2371_ _2361_ _2372_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4488__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3314__I _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__B1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4346__S _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6401__A2 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__I _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5912__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5704__I _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4748__C _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3454__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4810_ _1725_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6471__S _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _2342_ _2597_ _2603_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ mod.ldr_hzd\[4\] _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _1243_ _1476_ _1412_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6411_ _2356_ _3042_ _3047_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4706__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3623_ mod.registers.r8\[3\] _0416_ _0420_ mod.registers.r11\[3\] _0651_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6342_ _2999_ _3004_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3554_ _3170_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6273_ _0878_ _2893_ _2956_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3485_ _0508_ _0510_ _0511_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5614__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5224_ mod.pc_2\[13\] _2108_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout89_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _2140_ _2157_ _2158_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3693__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4106_ _0749_ _0750_ _0751_ _0752_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5086_ mod.rd_3\[1\] _2083_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4037_ mod.registers.r8\[14\] _0813_ _0898_ mod.registers.r6\[14\] _0893_ mod.registers.r12\[14\]
+ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_72_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _2722_ _2729_ _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4939_ _1844_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3748__A3 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _0242_ net55 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5524__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4308__S1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4633__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5189__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A3 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6090__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5361__A2 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3372__A1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3270_ _3118_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3675__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4494__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _2668_ mod.pc0\[5\] _2673_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6891_ _0118_ net200 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ mod.registers.r14\[7\] _2632_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4927__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5773_ _2507_ _2589_ _2592_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6129__A1 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _0711_ _0933_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4655_ _1110_ _1202_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3606_ _3175_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5352__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4586_ _1373_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6325_ _2659_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3537_ _0562_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5344__I _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6256_ _0591_ _2940_ _2945_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3468_ _0489_ _0492_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_103_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__S _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5207_ _2177_ _2034_ _2196_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6187_ _2899_ _2901_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3666__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3399_ _3211_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _2129_ _1914_ _2122_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3799__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5069_ net11 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3657__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__C1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__I _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4333__I _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6819__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout139_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _1216_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4371_ _1177_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5164__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A3 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3896__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _2830_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ _3149_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _2661_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3253_ mod.instr_2\[1\] _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__I mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6874_ _0101_ net205 mod.des.des_dout\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3820__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5825_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6499__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5756_ mod.registers.r12\[7\] _2578_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ mod.pc_2\[0\] _0527_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ mod.registers.r10\[14\] _2535_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _1663_ _1664_ _1665_ _1542_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4569_ _1110_ _1454_ _1209_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3887__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6308_ _2970_ _2977_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ mod.funct7\[2\] _2931_ _2903_ mod.instr\[20\] _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5802__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4836__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3639__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3750__C _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__B2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3575__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4772__B1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__A2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3590__A4 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3327__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4529__S _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_320 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_331 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_342 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_353 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_364 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6641__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3940_ _0578_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ mod.registers.r6\[11\] _0898_ _0817_ mod.registers.r13\[11\] _0899_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5610_ _2483_ _2484_ _2486_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6590_ _0223_ net92 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5555__A2 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3566__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _2382_ _2435_ _2439_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5472_ _2390_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4423_ _1125_ _1450_ _1402_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3407__I _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4354_ _1377_ _1378_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4381__I3 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ mod.instr_2\[10\] _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4285_ _1180_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5622__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__B2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout71_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _1891_ _2044_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_3236_ mod.des.des_counter\[1\] _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6283__A3 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6857_ _0084_ net135 mod.registers.r15\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5069__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout57 net61 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5808_ _2367_ _2610_ _2614_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout68 net86 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout79 net80 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _0015_ net172 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5739_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3745__C _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4506__B1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__B _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6514__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4285__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3493__B1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4592__B _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A1 _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _1095_ _1096_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4276__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__S _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4028__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4972_ _1932_ _1991_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5776__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _0344_ net76 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3923_ _0941_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6642_ _0275_ net64 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ mod.registers.r3\[11\] _0782_ _0800_ mod.registers.r6\[11\] _0882_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5528__A2 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3539__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _0206_ net89 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4736__C2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3785_ _0490_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5617__I _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _2415_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6537__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4406_ _0958_ _0729_ _0733_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5386_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5700__A2 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout203 net204 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3711__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _1359_ _1364_ _1257_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6687__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4268_ _1291_ _0942_ _0949_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_86_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5464__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ mod.pc\[9\] _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4199_ _1108_ _1218_ _1224_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4019__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5216__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3600__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5767__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6192__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__B _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5262__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6093__I _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__I _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout121_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3570_ _0597_ _0449_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3941__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3941__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__S _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5240_ _1106_ _2162_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ mod.des.des_dout\[28\] _2141_ _2170_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5172__I _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _0543_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4053_ _1080_ _1075_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 io_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3457__B1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__C _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _1932_ _1967_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__S _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _0933_ _0439_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _0258_ net66 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3837_ _3225_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4185__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _0189_ net120 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3768_ _0469_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3393__C1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _2329_ _2416_ _2419_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _3091_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3699_ _0706_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ mod.registers.r5\[11\] _2362_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5685__A1 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__I _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5369_ mod.registers.r4\[10\] _2317_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3448__B1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5988__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__B2 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4660__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4426__I _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6702__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6852__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5912__A2 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4723__I0 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4110__B _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4100__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout169_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ mod.ldr_hzd\[6\] _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ _1291_ _1320_ _1698_ _1164_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4167__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ mod.registers.r15\[7\] _3043_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3622_ mod.registers.r9\[3\] _0425_ _0429_ mod.registers.r10\[3\] _0650_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5903__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3914__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6341_ _1763_ _3000_ _3001_ _2983_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3553_ _3150_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ mod.pc_1\[11\] _2665_ _2955_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3484_ mod.registers.r11\[5\] _3164_ _0435_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5667__A1 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _2211_ _2217_ _2219_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3415__I _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ mod.registers.r1\[5\] _2146_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__I0 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ mod.pc_2\[0\] _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_56_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ _2092_ _1740_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4674__C _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _1060_ _1061_ _1062_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4690__B _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6395__A2 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5987_ _1926_ _2735_ _1941_ _1944_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6875__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4938_ _1837_ _1839_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4869_ _3101_ _1886_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5077__I _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6608_ _0241_ net91 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6539_ _0172_ net115 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__A1 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4881__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4156__I _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6138__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__I _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3235__I mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6748__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3675__A3 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6074__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5821__A1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4066__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _2682_ _2685_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6482__S _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _0117_ net198 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3832__B1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _2353_ _2631_ _2635_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4388__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ mod.registers.r12\[13\] _2590_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4723_ _1745_ _1746_ _1747_ _1748_ _1749_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4654_ _1678_ _1680_ _1681_ _1331_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3605_ mod.registers.r7\[2\] _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4585_ _0875_ _0951_ _3193_ _0837_ _1207_ _1269_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3899__B1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5625__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _2909_ _2977_ _2978_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3536_ _0540_ _0563_ _0443_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6255_ mod.pc_1\[5\] _2941_ _2942_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3467_ mod.registers.r10\[6\] _0493_ _0494_ mod.registers.r7\[6\] _0495_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4312__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ mod.pc_2\[11\] _2108_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6186_ _1860_ _2900_ _2891_ mod.instr\[1\] _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3398_ mod.registers.r5\[7\] _0423_ _0425_ mod.registers.r9\[7\] _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5137_ _1918_ _2120_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _2078_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4615__A2 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _1011_ _1046_ _1038_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3823__B1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4000__B1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5535__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4551__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4551__B2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4067__B1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4067__C2 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3814__B1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout201_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _1303_ _1395_ _1396_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__CLK net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3321_ _3141_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _2069_ _2763_ _2791_ _2792_ _2741_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_98_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ _3104_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6047__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4058__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6873_ _0100_ net208 mod.des.des_dout\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _2622_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5755_ _2489_ _2577_ _2581_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ mod.pc_2\[0\] _0527_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5686_ _2507_ _2534_ _2537_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ _1198_ _1212_ _1367_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4399__C _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _1373_ _1500_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__S _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3519_ _0428_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6307_ _2978_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1275_ _1250_ _1371_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6238_ _2930_ _2934_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4836__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ mod.instr\[20\] _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3759__B _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__A1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6277__A1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_310 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_321 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6029__A1 _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_332 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_343 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_354 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_365 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout151_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _0491_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6201__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3566__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ mod.registers.r7\[14\] _2436_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _2388_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5175__I _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4422_ _1428_ _1449_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4353_ _1248_ _1237_ _1241_ _1192_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3304_ mod.instr_2\[11\] _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_99_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4284_ _1215_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4818__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6023_ _2777_ _1891_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3235_ mod.des.des_counter\[0\] _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6283__A4 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6035__A4 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _0083_ net134 mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout58 net61 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5807_ mod.registers.r13\[10\] _2611_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3999_ mod.registers.r1\[12\] _0824_ _0992_ mod.registers.r13\[12\] _1027_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6787_ _0014_ net172 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4754__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ _2568_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ mod.registers.r10\[7\] _2523_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__B2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3493__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3493__B2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4164__I _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4993__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5170__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3720__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout199_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__B _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3484__A1 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A2 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _0779_ _1987_ _1990_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_51_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _0343_ net75 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3922_ _0948_ _0832_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4984__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _0274_ net53 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ mod.registers.r14\[11\] _0796_ _0454_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3539__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ mod.registers.r15\[8\] _0810_ _0811_ mod.registers.r3\[8\] _0812_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4736__B2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6572_ _0205_ net120 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5523_ _2357_ _2423_ _2428_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _2236_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _1188_ _0733_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5161__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _2100_ _2299_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4336_ _1210_ _1362_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xfanout204 net214 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3711__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout215 net1 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4267_ _1292_ _1294_ _0877_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6006_ _2704_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5464__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4198_ _1112_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4693__B _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__I _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4019__A3 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _0066_ net191 mod.ldr_hzd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4712__I _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3328__I _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6631__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6781__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4663__B1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5207__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5391__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout114_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3941__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _2152_ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4121_ _0521_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4052_ _1058_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3457__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput4 io_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _1900_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6504__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6159__B1 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3905_ _0635_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4885_ _1837_ _1839_ mod.pc\[3\] _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5628__I _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _0257_ net110 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3836_ mod.registers.r6\[9\] _0816_ _0863_ mod.registers.r1\[9\] _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5382__A1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4185__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3767_ mod.registers.r4\[8\] _0570_ _0794_ mod.registers.r1\[8\] _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6555_ _0188_ net120 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6654__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3393__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3393__C2 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5506_ mod.registers.r7\[0\] _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3698_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6486_ mod.des.des_dout\[36\] net8 _3078_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3592__B _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5437_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5363__I _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5685__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _2194_ _2316_ _2319_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4319_ _1333_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5299_ mod.registers.r3\[0\] _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3448__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3448__B2 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3611__I _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__I _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5273__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__I1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3687__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6476__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4100__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4670_ _1291_ _1315_ _1218_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__B _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3621_ mod.registers.r5\[3\] _0423_ _3226_ mod.registers.r2\[3\] _0418_ mod.registers.r6\[3\]
+ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4167__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ _0574_ _0575_ _0577_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6340_ _2999_ _3003_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6271_ _2709_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5116__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5183__I _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3483_ mod.registers.r5\[5\] _0460_ _3160_ mod.registers.r10\[5\] _0511_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ mod.registers.r1\[12\] _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3678__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5153_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4104_ _0748_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5084_ net12 _1828_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4035_ mod.registers.r10\[14\] _0991_ _0824_ mod.registers.r1\[14\] _1063_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4690__C _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5986_ mod.pc\[6\] _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ _1879_ _1957_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3602__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4262__I _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ mod.pc0\[2\] _1887_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5355__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _0240_ net94 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3819_ _0661_ _0845_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4799_ _1744_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6538_ _0171_ net117 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ mod.des.des_dout\[28\] net18 _3079_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3669__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3341__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4397__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3372__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A2 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout181_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3251__I mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3832__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__B _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3832__B2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ mod.registers.r14\[6\] _2632_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5585__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4388__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _2503_ _2589_ _2591_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4082__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4722_ _0714_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4653_ _1367_ _1482_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4810__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3604_ _3187_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4584_ _1526_ _1557_ _1270_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3899__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3899__B2 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6323_ _1765_ _2988_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3535_ mod.funct7\[0\] _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3426__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _0568_ _2940_ _2944_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3466_ _0430_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4848__B1 _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5205_ _2176_ _2202_ _2203_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6185_ _2896_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3397_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _2104_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6065__A2 _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _1713_ net22 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4076__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6842__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4018_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5576__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2722_ _2724_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__I0 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5879__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__B2 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5500__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4067__B2 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3814__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3814__B2 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__B1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6359__A3 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3290__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3578__B1 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5319__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6715__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3320_ mod.registers.r3\[7\] _3171_ _3172_ mod.registers.r6\[7\] _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3251_ mod.valid2 _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6865__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__B1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4077__I _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__B2 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _0099_ net208 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5823_ _2623_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5558__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3569__B1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5754_ mod.registers.r12\[6\] _2578_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4230__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4705_ _1729_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5636__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ mod.registers.r10\[13\] _2535_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _1325_ _1613_ _1186_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4533__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5730__A1 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _1373_ _1501_ _1228_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3741__B1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6306_ _1809_ _2965_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3518_ _3198_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _1460_ _1272_ _1335_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A2 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ mod.funct7\[1\] _2931_ _2903_ mod.instr\[19\] _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3449_ _3225_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _2885_ _2826_ _2886_ _2879_ _2880_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _2825_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5797__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3272__A2 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__S _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6738__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4772__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3980__B1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6277__A2 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4288__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_300 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_311 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_322 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_333 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_344 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_355 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_366 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__B _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4625__I _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4460__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout144_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5960__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3971__B1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5470_ _2343_ _2389_ _2395_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4421_ _1447_ _1146_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5712__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3723__B1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4352_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6268__A2 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3303_ _3141_ _3155_ _3133_ _3135_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4283_ mod.funct3\[0\] _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4279__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6022_ mod.pc\[11\] _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout57_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _0082_ net134 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5806_ _2364_ _2610_ _2613_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout59 net61 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6786_ _0013_ net170 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3998_ mod.registers.r9\[12\] _0805_ _0987_ mod.registers.r7\[12\] _0821_ mod.registers.r14\[12\]
+ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_5737_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4754__A2 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3962__B1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _2489_ _2522_ _2526_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4619_ _1239_ _1046_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4506__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5599_ _2477_ _2473_ _2478_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5219__B1 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4690__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3493__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5942__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4180__I _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4970_ _1988_ _1973_ _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _0854_ _0868_ _0872_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4984__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _0273_ net112 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3852_ mod.registers.r13\[11\] _0784_ _0788_ mod.registers.r15\[11\] _0880_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6186__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__B2 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4736__A2 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _0204_ net120 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3783_ _0478_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5522_ mod.registers.r7\[7\] _2424_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _2382_ _2375_ _2383_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4404_ _1429_ _1430_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5384_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout205 net206 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4335_ _1200_ _1289_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4266_ _0605_ _0778_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6005_ _1982_ _2719_ _2762_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4672__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4197_ _1220_ _3123_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4424__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4975__A2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6838_ _0065_ net183 mod.ldr_hzd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5924__A1 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _0399_ net174 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__I _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3519__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout107_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3254__I _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4120_ _0602_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4051_ _1042_ _1048_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_84_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3457__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 io_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__I _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _0596_ _1970_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3904_ _0454_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4884_ _1834_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6623_ _0256_ net107 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3835_ _3230_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3429__I _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6554_ _0187_ net122 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3766_ _3144_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3873__B _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3393__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5505_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3393__B2 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6485_ _3090_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3697_ _0707_ _0455_ _0719_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_106_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _2208_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5134__A2 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5367_ mod.registers.r4\[9\] _2317_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4318_ _1334_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5298_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4249_ _1274_ _1276_ _1270_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3448__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4723__I2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3687__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5061__A1 _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _0646_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4021__C1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__A3 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3551_ mod.registers.r10\[4\] _0578_ _0435_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _0911_ _2947_ _2954_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5116__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6313__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3482_ mod.registers.r13\[5\] _3140_ _0509_ mod.registers.r1\[5\] _0510_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5221_ _2117_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3678__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5152_ mod.des.des_dout\[26\] _2141_ _2151_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_69_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _0747_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6295__I _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4808__I _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5083_ mod.valid2 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4627__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4034_ mod.registers.r5\[14\] _0819_ _0823_ mod.registers.r2\[14\] _1062_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _2742_ _2706_ _2745_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5639__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ _1862_ _1951_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3602__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _1888_ _1889_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6606_ _0239_ net91 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3818_ mod.registers.r3\[9\] _0782_ _0797_ mod.registers.r10\[9\] _0846_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5355__A2 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4798_ _1773_ _1820_ _1821_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_20_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6771__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6537_ _0170_ net116 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5374__I _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3749_ _0775_ _0589_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__A1 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _3081_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5419_ _2356_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6399_ _2339_ _3035_ _3040_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3669__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4618__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5291__A1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5043__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5043__B2 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__S0 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6329__B _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4609__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout174_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A4 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3832__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ mod.registers.r12\[12\] _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _0710_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6794__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _1342_ _1679_ _1322_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6385__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3603_ mod.registers.r5\[2\] _0583_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4583_ _1349_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5194__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3899__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6322_ _2989_ _2990_ _2981_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3534_ _3198_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ mod.pc_1\[4\] _2941_ _2942_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3465_ _0428_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4848__A1 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ mod.registers.r1\[10\] _2185_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4848__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6184_ _2889_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout87_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _0412_ _3202_ _3204_ _3229_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_111_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5135_ _2102_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _2077_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4076__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4474__S _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4017_ _1044_ _0958_ _1023_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3823__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4273__I _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6222__B1 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _1908_ _1910_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4919_ _1836_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5899_ _2655_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6376__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3339__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4000__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3617__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4892__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3814__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5016__B2 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3578__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3527__I _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3750__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3250_ _3103_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4358__I _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3502__B2 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3262__I _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _0098_ net208 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4093__I _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5822_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3569__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5753_ _2487_ _2577_ _2580_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3569__B2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4230__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _1317_ _1721_ _1730_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4821__I _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _2503_ _2534_ _2536_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _1342_ _1336_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1358_ _1543_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5730__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3741__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _1796_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _0500_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3741__B2 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__I _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4497_ _1405_ _1444_ _1520_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6236_ _2930_ _2933_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3448_ mod.registers.r15\[6\] _0474_ _0475_ mod.registers.r12\[6\] _0476_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6167_ mod.des.des_dout\[19\] _2838_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3379_ _3203_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ mod.des.des_dout\[22\] _2105_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6098_ mod.instr\[2\] _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4049__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _2062_ _1074_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3980__A1 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3980__B2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__B1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3732__B2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5485__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_301 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_312 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_323 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_334 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_345 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5237__A1 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_356 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_367 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6393__I _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5737__I _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout137_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__B2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _1151_ _1152_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3723__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _1201_ _1281_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5472__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ _3154_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4282_ _1298_ _1299_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5476__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ _2770_ _2776_ _2660_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3487__B1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6009__S _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6854_ _0081_ net135 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ mod.registers.r13\[9\] _2611_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6785_ _0012_ net175 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6252__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ mod.registers.r10\[12\] _0991_ _0997_ mod.registers.r4\[12\] _0988_ mod.registers.r11\[12\]
+ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_22_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _2568_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3962__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5667_ mod.registers.r10\[6\] _2523_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3962__B2 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4618_ _0951_ _1616_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ mod.registers.r9\[1\] _2475_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4549_ _1273_ _1208_ _1474_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6219_ _2916_ _2922_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6705__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6855__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3705__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3705__B2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5292__I _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5458__A1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4130__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _0854_ _0873_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__B1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ mod.registers.r8\[11\] _0791_ _0797_ mod.registers.r10\[11\] _0879_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6186__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4197__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6570_ _0203_ net130 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3782_ _0474_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4304__C _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _2354_ _2423_ _2427_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ mod.registers.r5\[14\] _2376_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5697__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _1184_ _1263_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5383_ _2115_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4334_ _1093_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout206 net207 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5449__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4265_ _0840_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6004_ _2705_ _2761_ _2751_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4196_ _1111_ _1223_ _3131_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6728__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3450__I _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6878__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _0064_ net183 mod.ldr_hzd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6177__A2 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4281__I _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6768_ _0398_ net174 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5719_ _2497_ _2555_ _2558_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6699_ _0332_ net125 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6101__A2 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5860__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__I _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3871__B1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5612__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__B1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3474__I0 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A2 _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5679__A1 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3535__I mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4050_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5851__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4406__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _1971_ _1956_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3614__B1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3903_ _0546_ _0926_ _0930_ _0497_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6159__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ _3105_ _1726_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3834_ mod.registers.r13\[9\] _0817_ _0808_ mod.registers.r11\[9\] _0862_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6622_ _0255_ net108 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5906__A2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3917__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _0186_ net122 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3765_ mod.registers.r8\[8\] _0791_ _0792_ mod.registers.r2\[8\] _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5504_ _2414_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3393__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ mod.des.des_dout\[35\] net7 _3078_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3696_ _0720_ _0721_ _0722_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5435_ _2368_ _2361_ _2369_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4342__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _2184_ _2316_ _2318_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4317_ _1322_ _1341_ _1343_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _2271_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4248_ _0599_ _1266_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3908__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5835__I _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4723__I3 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5570__I _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5833__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3974__B _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4021__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4021__C2 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3550_ _3159_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6573__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3265__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3481_ _3143_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6313__A2 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4324__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5151_ _2152_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6077__A1 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4102_ _0703_ _0705_ _0725_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_57_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ net12 _2082_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4096__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ mod.registers.r9\[14\] _0805_ _0987_ mod.registers.r7\[14\] _1061_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4824__I _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6017__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2707_ _2744_ _2711_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5052__A2 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _0453_ _1953_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_21_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4260__B1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3602__A3 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4866_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _0238_ net104 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3817_ mod.registers.r8\[9\] _0791_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4797_ _1822_ _1823_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6536_ _0169_ net70 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3748_ _0763_ _0566_ _0588_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_106_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ mod.pc_2\[1\] _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6467_ mod.des.des_dout\[27\] net17 _3079_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4315__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _2173_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6398_ mod.registers.r15\[2\] _3037_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5349_ mod.registers.r4\[2\] _2305_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4618__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__S1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6596__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3357__A2 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6059__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5806__A1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout167_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5034__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4720_ mod.ldr_hzd\[15\] _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _1508_ _1646_ _1205_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3602_ _0623_ _0625_ _0627_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4545__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _1608_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4545__B2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3533_ _0554_ _0556_ _0557_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6321_ _2909_ _1812_ _2979_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6252_ _0676_ _2940_ _2943_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ mod.registers.r8\[6\] _0490_ _0491_ mod.registers.r6\[6\] _0420_ mod.registers.r11\[6\]
+ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_5203_ _2201_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4848__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ _2652_ _2898_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3395_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ _2103_ _2138_ _2139_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _1860_ _1740_ _1830_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_85_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ mod.pc_2\[12\] _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__B2 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ _2722_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4918_ _1855_ _1726_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5898_ _2675_ _1886_ _1894_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ mod.des.des_counter\[0\] _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4536__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3339__A2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6519_ _0152_ net42 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6289__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5053__C _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5264__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3275__A1 _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__A2 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__A1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__B2 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3578__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4775__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3750__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3543__I _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3502__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4374__I _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__D _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6870_ _0097_ net209 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ _2241_ _2567_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3569__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ mod.registers.r12\[5\] _2578_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4230__A3 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ _1653_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ mod.registers.r10\[12\] _2535_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4518__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4634_ _1302_ _1661_ _3132_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4565_ _1519_ _1349_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5191__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6304_ _1754_ _2974_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3516_ _0521_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3741__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4496_ _1125_ _1523_ _1401_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3447_ _3210_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6235_ mod.funct7\[0\] _2931_ _2927_ mod.instr\[18\] _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3453__I _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__B _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3378_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6166_ mod.instr\[19\] _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _2121_ _1859_ _2122_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6097_ _2832_ _2664_ _2833_ _2829_ _2831_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_111_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4049__A3 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5048_ _2062_ _1074_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__A1 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4233__B _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3980__A2 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6634__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5999__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_302 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_313 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_324 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_335 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_346 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_357 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_368 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3248__A1 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4194__I _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4922__I _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3420__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5173__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3474__S _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4350_ _1276_ _1251_ _1371_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3723__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3301_ mod.instr_2\[12\] _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _1286_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3273__I _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5476__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _2772_ _2773_ _2775_ _2757_ _2713_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3487__B2 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6425__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5228__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3239__A1 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4987__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6507__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _0080_ net211 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5928__I _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5804_ _2359_ _2610_ _2612_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout39 net40 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6784_ _0011_ net160 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _1012_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5735_ _2300_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6657__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _2487_ _2522_ _2525_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4617_ _1165_ _1414_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5597_ _2126_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _1415_ _1541_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4500__C _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4479_ _1460_ _1272_ _1207_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _0933_ _2917_ _2920_ mod.instr\[12\] _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6149_ mod.des.des_dout\[14\] _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6416__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__C _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3402__A1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5155__A1 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3705__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4130__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6407__A1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4138__B _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5748__I _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3850_ mod.pc_2\[11\] _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_32_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A2 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3781_ mod.registers.r10\[8\] _0547_ _0808_ mod.registers.r11\[8\] _0809_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5394__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5520_ mod.registers.r7\[6\] _2424_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5451_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4402_ _1139_ _1140_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_126_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ _2237_ _2322_ _2327_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4320__C _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__I _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4333_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout207 net210 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ _0832_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _2756_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4195_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout62_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3880__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__B _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__B _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3632__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6836_ _0063_ net172 mod.ldr_hzd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _0397_ net173 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3979_ _0985_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5718_ mod.registers.r11\[9\] _2556_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6698_ _0331_ net126 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5649_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5393__I _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3699__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3320__B1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3871__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3871__B2 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6822__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__B2 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3474__I1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5128__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__B1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4351__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4639__B1 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5300__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout197_I mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 io_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3862__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4951_ _0452_ _1953_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3614__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3614__B2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3902_ _0927_ _0928_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4882_ _1900_ _1896_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4315__C _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _0254_ net108 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5367__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3833_ _0856_ _0857_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3917__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6552_ _0185_ net72 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3764_ _3181_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5503_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4331__B _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _3089_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3695_ mod.registers.r7\[1\] _0632_ _0583_ mod.registers.r5\[1\] _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5434_ mod.registers.r5\[10\] _2362_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5365_ mod.registers.r4\[8\] _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5941__I _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4316_ _1203_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6258__B _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5296_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4247_ _1082_ _1231_ _0597_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6845__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4178_ _0569_ _1195_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3853__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3605__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4292__I _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _0046_ net180 mod.ri_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5358__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3908__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5530__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__I _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3844__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4416__B _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5298__I _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A3 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4021__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4021__B2 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6718__CLK net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout112_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3480_ mod.registers.r8\[5\] _0457_ _3152_ mod.registers.r9\[5\] _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5521__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__B1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _0527_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4377__I _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4101_ _0598_ _0602_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5081_ _2085_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4088__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4032_ mod.registers.r13\[14\] _0992_ _0997_ mod.registers.r4\[14\] _1060_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5983_ _2737_ _2743_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__B1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4934_ _0506_ _1934_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4260__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5001__I mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4865_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6001__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6604_ _0237_ net121 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3816_ _0842_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4012__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1756_ _1755_ _1754_ _1753_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6535_ _0168_ net42 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5760__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3747_ _0545_ _0566_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3456__I _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6466_ _3080_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3678_ _0703_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4315__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _2354_ _2347_ _2355_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5512__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__I _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _2336_ _3035_ _3039_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _2127_ _2303_ _2307_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__I _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5279_ _2202_ _2257_ _2261_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4079__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4787__C1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4750__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A1 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3366__I _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__A2 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3315__B _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3817__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _1237_ _1648_ _1677_ _1193_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput10 io_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3601_ mod.registers.r4\[2\] _0628_ _0499_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5742__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _1581_ _0644_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6690__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6320_ _1769_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3532_ mod.registers.r15\[4\] _0558_ _0559_ mod.registers.r5\[4\] _0560_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6298__A2 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6251_ mod.pc_1\[3\] _2941_ _2942_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5491__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3463_ _0417_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5202_ mod.des.des_dout\[31\] _2187_ _2198_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__3505__B1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6182_ _3114_ _2897_ _2891_ mod.instr\[0\] _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_97_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3394_ _3201_ _3217_ _3204_ _3228_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ mod.registers.r1\[3\] _2118_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5064_ _2059_ _1720_ _2074_ _2076_ _1103_ net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _1009_ _1006_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _1886_ _2723_ _1908_ _1910_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4917_ _1932_ _1933_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5897_ _2667_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3992__B1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4848_ _3102_ _1871_ _1872_ _1852_ _1874_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_20_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4536__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ mod.ldr_hzd\[6\] _1801_ _1803_ mod.ldr_hzd\[4\] _1798_ mod.ldr_hzd\[7\] _1807_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6518_ _0151_ net69 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ mod.des.des_dout\[20\] net5 _3066_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3275__A2 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6165__C _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6563__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4224__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5972__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4775__A2 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5820_ _2384_ _2616_ _2621_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _2483_ _2577_ _2579_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4702_ _1317_ _1720_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5682_ _2516_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4633_ _1654_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _1441_ _1432_ _1437_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6303_ _2975_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3515_ _0522_ _0527_ _0537_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_116_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4495_ _1493_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__I _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout92_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6234_ _2930_ _2932_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6140__A1 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3446_ _3206_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6165_ _2883_ _2875_ _2884_ _2879_ _2880_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3377_ _3204_ _3229_ _3222_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0730_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6586__CLK net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6096_ mod.des.des_dout\[1\] _2826_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _1044_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__C1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5949_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4757__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__I _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__B1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5706__A1 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3717__B1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4693__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_303 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_314 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_325 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_336 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_347 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_358 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_369 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3248__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4445__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4748__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3420__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3708__B1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5173__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3554__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3300_ mod.registers.r8\[7\] _3150_ _3152_ mod.registers.r9\[7\] _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _1302_ _1307_ _3132_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3487__A2 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3239__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _0079_ net209 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6189__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5803_ mod.registers.r13\[8\] _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5936__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ _0010_ net160 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3995_ _1017_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _2298_ _2441_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ mod.registers.r10\[5\] _2523_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5944__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _1342_ _1509_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _2470_ _2473_ _2476_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _1323_ _1458_ _1464_ _1340_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6113__A1 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4478_ _1407_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6217_ _2916_ _2921_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ _3150_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6148_ _2662_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6416__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6079_ _2794_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4427__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6015__I _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3402__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5854__I _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__C _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3780_ _0419_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5394__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _2230_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5146__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__B2 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _1190_ _0769_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5381_ mod.registers.r4\[15\] _2323_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4332_ _0729_ _0765_ _0958_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net210 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ _0938_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__B2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _2759_ _1994_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4194_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4329__B _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3880__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout55_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5939__I _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6624__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3632__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _0062_ net171 mod.ldr_hzd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3459__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6766_ _0396_ net173 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3978_ _1002_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6774__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5717_ _2493_ _2555_ _2557_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6697_ _0330_ net126 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5648_ _2241_ _2442_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5579_ _2444_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3699__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4896__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3320__B2 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3871__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3623__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3387__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5128__A2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4887__A1 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4887__B2 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5300__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__B2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _0452_ _1953_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3614__A2 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3901_ mod.registers.r2\[10\] _0865_ _0855_ mod.registers.r9\[10\] mod.registers.r14\[10\]
+ _0481_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__3279__I _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ _1736_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6620_ _0253_ net133 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3832_ mod.registers.r8\[9\] _0858_ _0859_ mod.registers.r3\[9\] _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6551_ _0184_ net73 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3763_ _0457_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6482_ mod.des.des_dout\[34\] net6 _3078_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3694_ mod.registers.r9\[1\] _0639_ _0578_ mod.registers.r10\[1\] _0722_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5433_ _2367_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4878__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5364_ _2304_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _1244_ _1239_ _1342_ _1199_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4246_ _1272_ _1273_ _1238_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3838__C1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4350__I0 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4177_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3853__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5055__A1 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__A1 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5358__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _0045_ net160 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _0379_ net188 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4030__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5530__A2 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__C _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3829__C1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3844__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__I _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3601__B _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5349__A2 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4021__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3827__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout105_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3532__B2 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _1007_ _1126_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5080_ _2086_ _2087_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5285__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4088__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ _1941_ _1944_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1954_ _1937_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4864_ _1842_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ mod.registers.r1\[9\] _0794_ _0792_ mod.registers.r2\[9\] _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6603_ _0236_ net121 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4342__B _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4795_ _1748_ _1747_ _1746_ _1745_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_119_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4012__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6534_ _0167_ net41 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3746_ _0598_ _0602_ _0544_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5760__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6465_ mod.des.des_dout\[26\] net16 _3079_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3677_ _0522_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6812__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ mod.registers.r5\[6\] _2348_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6396_ mod.registers.r15\[1\] _3037_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5512__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5347_ mod.registers.r4\[1\] _2305_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3472__I _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5278_ mod.registers.r2\[10\] _2258_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5276__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4079__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5901__B _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3826__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__B1 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__A1 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3514__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5267__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3817__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__B1 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4941__I _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A3 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3557__I _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3600_ _3176_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 io_in[1] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4580_ _1430_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5742__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3531_ _0422_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6250_ _2814_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3462_ _0415_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _2104_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3505__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3505__B2 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6181_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3393_ mod.registers.r8\[7\] _0416_ _0418_ mod.registers.r6\[7\] _0420_ mod.registers.r11\[7\]
+ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_69_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _2137_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _1848_ mod.des.des_counter\[1\] _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _0945_ _0956_ _1011_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_37_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ mod.pc\[3\] _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5430__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4916_ _1900_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5896_ _2669_ _1871_ _2674_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3992__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5168__B _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3992__B2 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _1873_ _1573_ _3098_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__A3 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4778_ mod.ldr_hzd\[5\] _1796_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3744__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6517_ _0150_ net69 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3729_ mod.registers.r13\[0\] _0576_ _0509_ mod.registers.r1\[0\] _0756_ _0757_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5682__I _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6448_ _3069_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5497__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4298__I _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6379_ mod.des.des_dout\[8\] net6 _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4247__B _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3680__B1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6858__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3983__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5592__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5488__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4999__B1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5412__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__I0 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5750_ mod.registers.r12\[4\] _2578_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4701_ _1309_ _1553_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3974__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5681_ _2514_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3287__I _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4632_ _1428_ _1449_ _0600_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4518__A3 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3726__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4563_ _1504_ _1580_ _1587_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4923__B1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3514_ _0539_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6302_ _1753_ _0003_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4494_ _1518_ _1447_ _0776_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5479__A1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6233_ _0657_ _2931_ _2927_ mod.instr\[17\] _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3445_ _0453_ _0456_ _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6164_ mod.des.des_dout\[18\] _2838_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3376_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _1861_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ mod.instr\[1\] _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1849_ _1001_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__B1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3662__C2 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5403__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6713__D _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5948_ _2697_ _1961_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__A1 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3965__B2 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5879_ _2654_ _2658_ _2660_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3717__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3717__B2 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6301__I _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4390__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4142__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6530__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4693__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_304 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_315 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_326 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_337 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_348 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_359 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6680__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3653__B1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3708__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3835__I _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__S _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4133__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4684__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3892__B1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5633__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6851_ _0078_ net211 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _2598_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ _1018_ _1019_ _1020_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6782_ _0009_ net161 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5733_ _2511_ _2561_ _2566_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _2483_ _2522_ _2524_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4615_ _1340_ _1479_ _1505_ _1325_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5595_ mod.registers.r9\[0\] _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4372__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4546_ _1553_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_2_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6553__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6113__A2 _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ _1439_ _0684_ _0643_ _0726_ _1206_ _1188_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4124__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3428_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6216_ _1750_ _2917_ _2920_ mod.instr\[11\] _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6147_ mod.instr\[14\] _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3359_ _3211_ _3205_ _3207_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4509__C _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6078_ _2777_ _2811_ _2818_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4427__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5624__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5029_ _1875_ _3094_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3635__B1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3938__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4060__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3402__A3 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5870__I _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4115__A1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5863__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3390__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A2 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A1 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout135_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4729__I0 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _1148_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5380_ _2231_ _2322_ _2326_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _1356_ _1357_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5780__I _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4106__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout209 net210 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4262_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4657__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ mod.pc\[8\] _1857_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ mod.funct3\[1\] _3122_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_67_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4409__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3632__A3 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _0061_ net170 mod.ldr_hzd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5020__I _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A1 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _0395_ net173 mod.instr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3977_ _1003_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5955__I _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4593__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ mod.registers.r11\[8\] _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _0329_ net76 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _2511_ _2504_ _2512_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _2371_ _2458_ _2463_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4896__A2 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5904__B _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4529_ _1439_ _0684_ _1335_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A2 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3856__B1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3320__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6599__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4033__B1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4336__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4639__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 io_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_64_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ mod.registers.r1\[10\] _0863_ _0808_ mod.registers.r11\[10\] _0928_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4880_ _0676_ _1901_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_60_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _3223_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ _0183_ net71 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3762_ _0783_ _0785_ _0787_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__3509__B _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5501_ _2270_ _2299_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _3088_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3693_ mod.registers.r14\[1\] _0624_ _0626_ mod.registers.r11\[1\] _0721_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _2201_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5363_ _2302_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ _1326_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _2090_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5827__A1 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ _0589_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3838__B1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3838__C2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4176_ _0706_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__I _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5055__A2 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6252__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6741__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _0044_ net161 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4566__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6748_ _0378_ net187 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ _0312_ net82 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4869__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5818__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3829__B1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3829__C2 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A2 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6614__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3532__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5809__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _1052_ _1057_ _0834_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6764__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__C _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ mod.pc\[5\] _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4932_ _0506_ _1934_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3599__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__A1 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4863_ _1833_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4548__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ _0235_ net131 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3814_ mod.registers.r14\[9\] _0796_ _0800_ mod.registers.r6\[9\] _0842_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4794_ _1761_ _1763_ _1758_ _1781_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_6533_ _0166_ net71 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3745_ _0727_ _0762_ _0772_ _0682_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3676_ _3106_ _0502_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4849__I mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5415_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6395_ _2328_ _3035_ _3038_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3753__I _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5346_ _2116_ _2303_ _2306_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _2194_ _2257_ _2260_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4228_ _1201_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ _0932_ _0729_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6637__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5267__A2 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__B2 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__B _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A4 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput12 io_in[2] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout215_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3530_ _3206_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3461_ mod.registers.r5\[6\] _0487_ _0488_ mod.registers.r9\[6\] _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5200_ _1934_ _2153_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3505__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6180_ _2793_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3392_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5131_ mod.des.des_dout\[24\] _2105_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _2073_ _2074_ _2075_ net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4013_ _1039_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A1 _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6207__B2 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5966__B1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5964_ _1888_ _2719_ _2726_ _2727_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _0506_ _1934_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_80_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5895_ _2670_ mod.pc0\[1\] _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _1858_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3992__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__I _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4777_ mod.ldr_hzd\[2\] _1802_ _1803_ mod.ldr_hzd\[0\] _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6516_ _0149_ net43 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3744__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3728_ _0742_ _0634_ _3188_ _0636_ _0743_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6447_ mod.des.des_dout\[19\] net4 _3066_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3659_ mod.registers.r1\[1\] _3231_ _3219_ mod.registers.r4\[1\] _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _3016_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3901__C1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5329_ mod.registers.r3\[12\] _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__A2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4457__B1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5203__I _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__B2 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__B1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__C1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__I0 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3983__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4932__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__I _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__B2 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3671__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout165_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6802__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3423__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3568__I mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4700_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3974__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _2501_ _2528_ _2533_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _1290_ _1656_ _1657_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3726__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _1289_ _1583_ _1589_ _3131_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6301_ _2973_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3513_ _3194_ _0540_ _0443_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4493_ _1444_ _1520_ _1120_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ _2796_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3444_ _0463_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ mod.instr\[18\] _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3375_ mod.instr_2\[14\] _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _2112_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6094_ _2824_ _2664_ _2827_ _2829_ _2831_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_fanout78_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__I mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _2059_ _1392_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3662__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__B2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__B _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5403__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5947_ _2703_ _2706_ _2712_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3414__A1 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3965__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5167__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ _1855_ _1829_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5693__I _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3717__A2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_305 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_316 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_327 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_338 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_349 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6825__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__I _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__B2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3388__I _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3708__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4947__I _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4684__A3 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3892__A1 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3892__B2 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5633__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3644__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__I _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__B _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6850_ _0077_ net209 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _2596_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6781_ _0008_ net182 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3993_ mod.registers.r5\[12\] _0967_ _0972_ mod.registers.r2\[12\] _1021_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5732_ mod.registers.r11\[15\] _2562_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5663_ mod.registers.r10\[4\] _2523_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__I _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _1344_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5594_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4545_ _1563_ _1569_ _1572_ _1400_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4372__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4476_ _1181_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6215_ _2890_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6848__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6146_ _2869_ _2863_ _2870_ _2867_ _2868_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ mod.instr_2\[15\] _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ mod.pc_1\[11\] _2812_ _2815_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3289_ _3141_ _3137_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__A3 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _2036_ _2044_ _2001_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input10_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__B _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3635__B2 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4060__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4363__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3571__B1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5312__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__A1 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3626__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3626__B2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4729__I1 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ _1190_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4106__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _1124_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _2753_ _2719_ _2758_ _2741_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_79_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6833_ _0060_ net171 mod.ldr_hzd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6764_ _0394_ net170 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4042__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3976_ _0427_ _0829_ _0902_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6520__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5715_ _2543_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5790__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6695_ _0328_ net76 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3756__I _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5646_ mod.registers.r9\[15\] _2505_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5542__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5577_ mod.registers.r8\[11\] _2459_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6670__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _1261_ _1267_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4459_ _1396_ _1486_ _1289_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3856__B2 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ mod.des.des_dout\[9\] _2848_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__B1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3608__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__A2 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5211__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4033__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4033__B2 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3387__A3 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6089__A2 _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4272__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6543__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3830_ _0415_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3761_ mod.registers.r7\[8\] _0585_ _0788_ mod.registers.r15\[8\] _0789_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5772__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6693__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ _2385_ _2408_ _2413_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ mod.des.des_dout\[33\] net5 _3084_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3692_ mod.registers.r15\[1\] _0518_ _0582_ mod.registers.r3\[1\] _0720_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _2365_ _2361_ _2366_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5791__I _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _2174_ _2310_ _2315_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _1323_ _1337_ _1340_ _1197_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _2269_ _2240_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4244_ _0593_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3838__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4175_ _1199_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6252__A2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _0043_ net147 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5763__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _0377_ net187 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3959_ _0494_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6678_ _0311_ net83 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4318__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ mod.registers.r9\[10\] _2495_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3526__B1 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3829__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6243__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__I _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5754__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__B1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5506__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout195_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5980_ _1927_ _2719_ _2740_ _2741_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4931_ _0903_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5993__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ mod.pc\[2\] _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6601_ _0234_ net123 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3813_ mod.pc_2\[9\] _0661_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5745__A1 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _1767_ _1768_ _1765_ _1769_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_119_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6532_ _0165_ net39 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3744_ _0770_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3675_ _0562_ _0689_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5414_ _2166_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ mod.registers.r15\[0\] _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5345_ mod.registers.r4\[0\] _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ mod.registers.r2\[9\] _2258_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6589__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4865__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4227_ _1193_ _1233_ _1237_ _1241_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_29_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4484__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4158_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4086__B _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4236__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4089_ _3120_ _3109_ _1116_ _3111_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4105__I mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3944__I _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4475__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4778__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__B1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__C _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput13 io_in[3] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4950__A2 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout110_I net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout208_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3460_ _0424_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6731__CLK net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4702__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3391_ _0413_ _0414_ _3221_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5130_ _0676_ _2107_ _2122_ _2135_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__I _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _0000_ _1851_ _1069_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4466__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6881__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ _1024_ _1038_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3513__I0 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5966__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _2650_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4634__B _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _1935_ _1922_ _1936_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5894_ _2080_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4353__C _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4845_ _0689_ _0702_ _1849_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3729__B1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4776_ mod.instr_2\[5\] _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6515_ _0148_ net42 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3727_ mod.registers.r5\[0\] _0583_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3764__I _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6446_ _3068_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3658_ _0644_ _0682_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6143__B2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6377_ _3026_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3589_ mod.registers.r13\[2\] _0480_ _0481_ mod.registers.r14\[2\] _0616_ _0617_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5328_ _2274_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3901__B1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3901__C2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__B _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4595__I _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _2133_ _2244_ _2249_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4457__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4457__B2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__A1 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5957__B2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3939__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__B1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__C2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4480__I1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3499__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4999__A2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout190 net194 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3671__A2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3423__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _1656_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4561_ _1124_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4923__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6300_ _2677_ _1744_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3512_ mod.funct7\[1\] _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4492_ _1493_ _1519_ _0590_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6231_ _2651_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3443_ _0465_ _0466_ _0468_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6162_ _2881_ _2875_ _2882_ _2879_ _2880_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ mod.registers.r4\[7\] _3219_ _3224_ mod.registers.r3\[7\] mod.registers.r2\[7\]
+ _3226_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_112_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4629__B _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5113_ _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6093_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5044_ _2021_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__I mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _2707_ _2708_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3414__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _2649_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _1836_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5167__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__I _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _1785_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6429_ _2381_ _3054_ _3058_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4678__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4539__B _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__I _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_306 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_317 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_328 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_339 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3653__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__I _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4602__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__B2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A3 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3892__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5800_ _2356_ _2604_ _2609_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6780_ _0007_ net167 mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ mod.registers.r8\[12\] _0971_ _0962_ mod.registers.r7\[12\] _1020_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _2509_ _2561_ _2565_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ _2516_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6346__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4613_ _1596_ _1640_ _1367_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5593_ _2471_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4203__I _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4544_ _1570_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1229_ _1502_ _1203_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ _2916_ _2919_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout90_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3426_ _3167_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3868__C1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3332__A1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ mod.des.des_dout\[13\] _2860_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3357_ _3208_ _3209_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _2019_ _2811_ _2817_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3288_ mod.instr_2\[13\] _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__A4 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _2037_ _2034_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_73_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3635__A2 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4094__B _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _2697_ _2045_ _2671_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4822__B _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6337__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6337__B2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4348__B1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3571__B2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5312__A2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3323__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5076__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3399__I _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__B _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6328__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4729__I2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5119__I _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5551__A2 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3562__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4958__I _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _3132_ _1122_ _1174_ _1283_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_99_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4106__A3 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4191_ _3120_ _3128_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4814__A1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _0059_ net192 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _0393_ net175 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3975_ _0932_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4042__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6413__I _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _2541_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _0327_ net74 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5790__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _2236_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5576_ _2368_ _2458_ _2462_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4527_ _1339_ _1526_ _1554_ _1209_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3772__I _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4458_ _0840_ _1154_ _1159_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4089__B _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3409_ _3110_ _3113_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4389_ _1119_ _1202_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_58_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3856__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6128_ mod.instr\[9\] _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5058__B2 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6059_ _1927_ _2803_ _2806_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3608__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3947__I _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4033__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6495__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A3 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3847__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5049__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__S _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4018__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3480__B1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout140_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6838__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3760_ _3185_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5772__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ _0708_ _0709_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5430_ mod.registers.r5\[9\] _2362_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5361_ mod.registers.r4\[7\] _2311_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _1339_ _1242_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5292_ _2099_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5288__A1 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _1262_ _1268_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3838__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _1200_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4637__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6815_ _0042_ net147 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4372__B _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _0376_ net186 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3958_ _0804_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5763__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6677_ _0310_ net83 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3889_ mod.registers.r9\[10\] _0781_ _0788_ mod.registers.r15\[10\] _0917_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _2201_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3526__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3526__B2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5559_ _2444_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__A1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3829__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4254__A2 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4282__B _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3765__A1 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__B2 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout188_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5132__I _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6660__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _0486_ _0496_ _1915_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4796__A3 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ _1834_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6600_ _0233_ net70 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3812_ _0832_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4792_ _1774_ _1792_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6531_ _0164_ net45 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3743_ _0619_ _0620_ _0642_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6462_ mod.des.des_counter\[2\] _2076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3674_ _0690_ _0691_ _0692_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _2351_ _2347_ _2352_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6393_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5307__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4211__I _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4308__I0 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5275_ _2184_ _2257_ _2259_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4226_ _1243_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4157_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3692__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4088_ mod.funct7\[1\] _3114_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4236__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5977__I _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3747__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6729_ _0359_ net141 mod.pc0\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4944__B1 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4121__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3960__I _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5887__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5975__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__B2 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput14 io_in[4] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4031__I _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout103_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3910__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3870__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _3097_ _3093_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4011_ _1024_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4466__A2 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6833__D _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _2705_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ _1918_ _1919_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5893_ _2669_ _1847_ _2672_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4206__I _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _1857_ _1866_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5718__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3729__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3729__B2 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _1793_ mod.instr_2\[3\] _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6514_ _0147_ net43 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3726_ mod.registers.r7\[0\] _0632_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4529__I0 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6445_ mod.des.des_dout\[18\] net3 _3066_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6143__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3657_ _0683_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6376_ mod.des.des_dout\[7\] net5 _3022_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3588_ _0612_ _3208_ _0613_ _0614_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3901__A1 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__I _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5327_ _2272_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3901__B2 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3780__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ mod.registers.r2\[2\] _2246_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5654__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4209_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5189_ _2177_ _1999_ _2149_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3968__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__B2 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4696__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout180 net181 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout191 net193 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A3 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5410__I _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A1 _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4620__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__B1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4470__B _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3865__I _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4560_ _0772_ _1138_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4491_ _0686_ _0773_ _1518_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4136__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3442_ mod.registers.r14\[6\] _0469_ _3185_ mod.registers.r15\[6\] _0470_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6230_ _2923_ _2929_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ mod.des.des_dout\[17\] _2872_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3373_ _3225_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__B1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _1861_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6092_ _2649_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A2 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1966_ _2048_ _2049_ _1851_ _2058_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6061__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4072__B1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _2657_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _3102_ _1847_ _1850_ _1852_ _1854_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__I mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4375__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _1746_ _1775_ _1778_ _1745_ _1779_ _1747_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ mod.registers.r1\[0\] _3231_ _3218_ mod.registers.r4\[0\] _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4689_ _1094_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6428_ mod.registers.r15\[14\] _3055_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4678__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3724__B _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6359_ _3092_ _3093_ mod.des.des_counter\[2\] _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3886__B1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5627__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_307 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_318 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_329 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6052__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6871__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4118__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5405__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5618__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5140__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ mod.registers.r13\[12\] _0959_ _0965_ mod.registers.r1\[12\] _1019_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ mod.registers.r11\[14\] _2562_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _2514_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _1092_ _1377_ _1363_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5592_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _1208_ _1118_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4109__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _1500_ _1501_ _0621_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5857__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _1749_ _2917_ _2913_ mod.instr\[10\] _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3425_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3868__B1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3868__C2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3332__A2 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6144_ mod.instr\[13\] _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout83_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3356_ _3203_ mod.instr_2\[14\] _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5609__A1 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ mod.pc_1\[10\] _2812_ _2815_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3287_ _3139_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _2037_ _2042_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4375__B _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6744__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4832__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ _2677_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _2378_ _2643_ _2646_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4348__A1 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3556__C1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5848__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3859__B1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4520__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3323__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3626__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4587__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4732__C _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6328__A2 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4729__I3 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6617__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3562__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__A1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5135__I _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6767__CLK net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A2 _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6831_ _0058_ net192 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4027__B1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__A1 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _0392_ net176 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3974_ _0986_ _1001_ _0827_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4642__C _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5713_ _2491_ _2549_ _2554_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6693_ _0326_ net76 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4214__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5644_ _2509_ _2504_ _2510_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5575_ mod.registers.r8\[10\] _2459_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4526_ _1355_ _1275_ _1250_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _1286_ _1446_ _1467_ _1469_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__4089__C _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4502__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3408_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4388_ _1414_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6127_ _2853_ _2851_ _2854_ _2855_ _2856_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ _3169_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5058__A2 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6255__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ mod.pc_1\[4\] _2805_ _2799_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _2007_ _2023_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__B _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__C _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5049__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3480__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3480__B2 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout133_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _3125_ _0713_ _0716_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4732__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _2167_ _2310_ _2314_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4311_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5291_ _2237_ _2263_ _2268_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4242_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _0683_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4209__I _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5996__B1 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout46_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _0041_ net147 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6745_ _0375_ net145 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3957_ _0957_ _0958_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _0309_ net59 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3888_ _0912_ _0913_ _0914_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5627_ _2497_ _2494_ _2498_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3783__I _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3526__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _2343_ _2445_ _2451_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4509_ _1521_ _1524_ _1525_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5489_ mod.registers.r6\[11\] _2403_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5503__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4119__I _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__B1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__C1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6334__I _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3765__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4738__B _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4457__C _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4796__A4 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4860_ _3105_ _1838_ _1885_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_33_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3811_ _0837_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4791_ _1810_ _1818_ _1774_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6530_ _0163_ net44 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3742_ _0763_ _0765_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4953__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _3076_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3673_ _0697_ _0698_ _0699_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4705__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ mod.registers.r5\[5\] _2348_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6392_ _3033_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _2301_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4308__I1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ mod.registers.r2\[8\] _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ _1244_ _1248_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5130__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3692__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3692__B2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ _1113_ _1079_ _1081_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_71_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__I _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4989_ _2005_ _2006_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6728_ _0358_ net148 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3747__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__B2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _0292_ net60 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput15 io_in[5] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3637__B _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__B _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5360__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4466__A3 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4010_ _0827_ _1033_ _1036_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_78_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4982__I _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _2722_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_92_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4474__I0 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3598__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__B1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4912_ _1918_ _1919_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_45_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__A2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _2670_ mod.pc0\[0\] _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _1867_ _1835_ _1845_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6513_ _0146_ net41 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3725_ _0749_ _0750_ _0751_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5318__I _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6444_ _3067_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4529__I1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3656_ _0680_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5351__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _3025_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3587_ mod.registers.r15\[2\] _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5326_ _2209_ _2286_ _2291_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3901__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5257_ _2127_ _2244_ _2248_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4208_ _1234_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _2005_ _2178_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _0874_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_44_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5002__B _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6500__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout170 net171 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout181 net185 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout192 net193 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6445__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3671__A4 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4307__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6070__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4243__S _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4908__B2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__B1 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5581__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout213_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3510_ _3107_ _3165_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4490_ _0777_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4136__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A1 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3441_ _3183_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6381__I0 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6160_ mod.instr\[17\] _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3372_ _3211_ _3220_ _3222_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__B2 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _2103_ _2116_ _2119_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _2828_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _3100_ _2054_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4217__I _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A2 _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5944_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4072__B2 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6523__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5875_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4826_ _1853_ _1733_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _1748_ _1777_ _0694_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3583__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3708_ mod.registers.r7\[0\] _0431_ _3224_ mod.registers.r3\[0\] _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4688_ _1105_ _1107_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6427_ _2378_ _3054_ _3057_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5324__A1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6372__I0 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3791__I _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3639_ mod.registers.r5\[3\] _0460_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6358_ _3014_ _3015_ _2727_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3886__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3886__B2 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ mod.registers.r3\[4\] _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6289_ _2965_ _2966_ _2895_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_308 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_319 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4127__I _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5563__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5315__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__I0 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__A2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout163_I net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ mod.registers.r15\[12\] _0981_ _0978_ mod.registers.r12\[12\] _1018_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _2481_ _2515_ _2521_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _1040_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5554__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5591_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _1435_ _1564_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4762__C1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4109__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5306__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _0875_ _1246_ _0837_ _0951_ _1338_ _1265_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6212_ _2916_ _2918_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3424_ mod.pc_2\[6\] _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3868__A1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6143_ _2865_ _2863_ _2866_ _2867_ _2868_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3355_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout76_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _2014_ _2811_ _2816_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3286_ _3134_ _3136_ _3138_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ _2039_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5085__A3 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5927_ _2670_ mod.pc0\[11\] _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4596__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5793__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ mod.registers.r14\[13\] _2644_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4348__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5545__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5789_ mod.registers.r13\[3\] _2599_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3556__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3556__C2 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3859__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3859__B2 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3470__B _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6273__A2 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5536__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6021__B _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _0057_ net192 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4027__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4027__B2 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6761_ _0391_ net175 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4578__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5775__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3973_ _0995_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_62_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3786__B1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5712_ mod.registers.r11\[7\] _2550_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6692_ _0325_ net53 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5643_ mod.registers.r9\[14\] _2505_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5527__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _2365_ _2458_ _2461_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4525_ _1401_ _1539_ _1549_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4456_ _1470_ _1471_ _1482_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6711__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3407_ _3166_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4387_ _1109_ _1355_ _1235_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _2830_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _3173_ _3182_ _3186_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_100_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6157__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4266__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3269_ mod.funct3\[0\] _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6861__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _2024_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3529__B1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5236__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6067__I _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4516__S _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4743__C _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3480__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5509__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4251__S _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6182__B2 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4310_ _1187_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5290_ mod.registers.r2\[15\] _2264_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ _0706_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4496__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4172_ _0567_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4248__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5996__A1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5996__B2 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6813_ _0040_ net157 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout39_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _0374_ net150 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3956_ _0970_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6675_ _0308_ net87 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4971__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3887_ mod.registers.r7\[10\] _0585_ _0677_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5626_ mod.registers.r9\[9\] _2495_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5557_ mod.registers.r8\[3\] _2447_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4508_ _1504_ _1532_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _2368_ _2402_ _2406_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4895__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _1457_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6109_ _2828_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5987__B2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__B1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6607__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3998__C2 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4135__I _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4478__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__C _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4754__B _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4246__S _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _0828_ _0831_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _1811_ _1813_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _0766_ _0661_ _0767_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__4953__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ mod.des.des_dout\[25\] net10 _3060_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3672_ mod.registers.r15\[1\] _3206_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5411_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _3034_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3913__B1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5342_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5273_ _2245_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4308__I2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4224_ _1244_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5130__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4155_ _1003_ _0660_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3692__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _1079_ _1081_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A1 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4988_ _2005_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6727_ _0357_ net144 mod.pc0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3939_ _0460_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6146__B2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _0291_ net59 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ mod.registers.r9\[4\] _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6589_ _0222_ net89 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__B _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3743__B _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3380__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5514__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3969__I _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6345__I _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A2 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__I _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 io_in[6] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__A1 _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5424__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6456__S _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout193_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _1886_ _2723_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4474__I1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4623__B2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4911_ _0935_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5891_ _2080_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ mod.pc\[1\] _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5179__A2 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4773_ _1797_ mod.instr_2\[3\] _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3724_ mod.registers.r4\[0\] _0628_ _0499_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6512_ _0145_ net95 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ mod.des.des_dout\[17\] net2 _3066_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3655_ _0456_ _0660_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6374_ mod.des.des_dout\[6\] net4 _3022_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5351__A2 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3586_ _3215_ _0414_ _3232_ _3205_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5325_ mod.registers.r3\[11\] _2287_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6300__A1 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ mod.registers.r2\[1\] _2246_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4207_ _1189_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _2087_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _1165_ _0873_ _0803_ _0838_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4394__B _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input19_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4069_ mod.registers.r9\[15\] _0805_ _0988_ mod.registers.r11\[15\] _1097_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4614__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4917__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4473__S0 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__B _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__A1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout160 net163 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout171 net172 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout182 net183 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout193 net194 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__I _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5030__B2 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3592__A1 _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout206_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3440_ mod.registers.r7\[6\] _0467_ _3189_ mod.registers.r12\[6\] _0468_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6381__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3371_ _3223_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5110_ mod.registers.r1\[0\] _2118_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ net13 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ mod.pc0\[12\] _1909_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4844__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3647__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5943_ _2079_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4072__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _2655_ _1828_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4825_ _1848_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5021__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6818__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _1776_ _1780_ _1782_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3583__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3707_ _0703_ _0705_ _0725_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3583__B2 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4687_ _3121_ _1712_ _1714_ _1317_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6426_ mod.registers.r15\[13\] _3055_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3638_ _0662_ _0663_ _0664_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6372__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3569_ _0596_ _0436_ _3169_ _3191_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6357_ _2908_ _2986_ _3008_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3886__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _2274_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6288_ mod.ins_ldr_3 _2936_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_309 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _2178_ _2059_ _1720_ _2163_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_76_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3513__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__B _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5260__A1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3810__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6498__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5012__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3574__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5315__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__B1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3877__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A1 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout156_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__B1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _1126_ _1320_ _1637_ _1319_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5590_ _2100_ _2442_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5554__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3565__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4541_ _1400_ _1565_ _1566_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__4762__B1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__C2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4472_ _1092_ _1058_ _1009_ _1024_ _1264_ _1204_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4109__A3 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5306__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3423_ _3193_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6211_ _1713_ _2917_ _2913_ mod.instr\[9\] _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3868__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6142_ _2830_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3354_ _3200_ mod.instr_2\[16\] _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ mod.pc_1\[9\] _2812_ _2815_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3285_ mod.instr_2\[13\] _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _0878_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4293__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__B _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4045__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6640__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ _2678_ _2031_ _2695_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5857_ _2373_ _2643_ _2645_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _3104_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5788_ _2339_ _2597_ _2602_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3556__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6790__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3556__B2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ mod.ldr_hzd\[7\] _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3308__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3308__B2 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _2353_ _3042_ _3046_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3307__I _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3859__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5233__A1 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5784__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3547__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3547__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4757__B _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4249__S _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__I _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6663__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4027__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A1 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6760_ _0390_ net175 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5775__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3972_ _0996_ _0998_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3786__A1 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ _2489_ _2549_ _2553_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3786__B2 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6691_ _0324_ net39 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5642_ _2230_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ mod.registers.r8\[9\] _2459_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5607__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _1483_ _1513_ _1551_ _1400_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _1454_ _1330_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3406_ _3199_ _0411_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4386_ _1335_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3710__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6125_ _2828_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ mod.registers.r7\[7\] _3187_ _3189_ mod.registers.r12\[7\] _3190_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5342__I _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3268_ _3120_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6056_ _2793_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4266__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6374__S _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _2007_ _2023_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A3 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ _2683_ mod.pc0\[4\] _2684_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6889_ _0116_ net199 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3529__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3529__B2 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6536__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6686__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5206__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5509__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6182__A2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4193__A1 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ _1263_ _1266_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4171_ _1092_ _1118_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__A2 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _0039_ net157 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3759__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6743_ _0373_ net144 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3955_ _0973_ _0976_ _0979_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6674_ _0307_ net60 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4971__A3 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3886_ mod.registers.r13\[10\] _0784_ _0794_ mod.registers.r1\[10\] _0914_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5625_ _2193_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5337__I _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4241__I _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5556_ _2340_ _2445_ _2450_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4507_ _1380_ _1374_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5487_ mod.registers.r6\[10\] _2403_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _1459_ _1462_ _1465_ _1257_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4369_ _1395_ _1396_ _1303_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3695__B1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6108_ mod.des.des_dout\[4\] _2835_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4239__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6484__I0 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _2788_ _2790_ _2739_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__B2 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4175__A1 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4478__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5427__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__B1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4754__C _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _0631_ _0633_ _0638_ _0640_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3610__B1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _0427_ _0695_ mod.registers.r13\[1\] _0694_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6851__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4166__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _2156_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3913__B2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5341_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5272_ _2243_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4308__I3 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5106__B _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ _0875_ _1245_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4085_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5620__I _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout51_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6394__A2 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _0441_ _1034_ _1035_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6451__I _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _0356_ net150 mod.pc0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3938_ mod.registers.r1\[13\] _0965_ _0436_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6146__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ _0290_ net54 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3869_ mod.registers.r1\[11\] _0863_ _0808_ mod.registers.r11\[11\] _0897_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ _2474_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6588_ _0221_ net130 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5539_ _2379_ _2435_ _2438_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4880__A2 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6724__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4632__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6874__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 io_in[7] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5896__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4699__A2 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__I _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5648__A1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3659__B1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4871__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3674__A3 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout186_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ _1858_ _1537_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5890_ _2667_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _1843_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6271__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4387__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4772_ mod.ldr_hzd\[1\] _1796_ _1799_ mod.ldr_hzd\[3\] _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6511_ _0144_ net87 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3723_ mod.registers.r11\[0\] _0626_ _0571_ mod.registers.r2\[0\] _0751_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6442_ _3060_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3654_ _0674_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _3024_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3585_ _3209_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4659__C _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ _2202_ _2286_ _2290_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout99_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5255_ _2116_ _2244_ _2247_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4206_ _0706_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _2176_ _2184_ _2186_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6747__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _0854_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__C _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ mod.registers.r13\[15\] _0992_ _0987_ mod.registers.r7\[15\] _0821_ mod.registers.r14\[15\]
+ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_43_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3822__B1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4378__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6181__I _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _0342_ net77 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5525__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3889__B1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4302__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout150 net154 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout161 net163 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout172 net177 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout183 net185 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout194 net195 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6091__I _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3416__I0 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3592__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout101_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3370_ _3221_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_124_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__S _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _2055_ _1928_ _1892_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4844__A2 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A1 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5942_ _1739_ _1840_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_46_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ net12 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5021__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ mod.ldr_hzd\[11\] _1777_ _1775_ mod.ldr_hzd\[9\] _1779_ mod.ldr_hzd\[10\]
+ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3706_ _0545_ _0729_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3583__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__A1 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _1713_ _1708_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6425_ _2373_ _3054_ _3056_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3637_ mod.registers.r4\[3\] _3177_ _3167_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4532__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ _1748_ _3006_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3568_ mod.pc_2\[7\] _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_115_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _2272_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6287_ _1774_ _2661_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3499_ _0439_ _0525_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _2211_ _2231_ _2232_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _1880_ _2153_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6037__A1 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3749__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A2 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3574__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3484__B _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4523__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__B2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6086__I mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4826__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__B1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6200__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _1130_ _1222_ _1567_ _0735_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3565__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__A1 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__B2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4471_ _1329_ _1395_ _1160_ _1468_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6210_ _2796_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4514__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3422_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6141_ net13 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3353_ _3201_ _3202_ _3204_ _3205_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3284_ mod.instr_2\[12\] _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _0563_ _1034_ _1035_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3413__I _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5242__A2 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4045__A3 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5925_ _2668_ mod.pc0\[10\] _2673_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4244__I _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ mod.registers.r14\[12\] _2644_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4807_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ mod.registers.r13\[2\] _2599_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3556__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ _1765_ _1759_ _0933_ _3147_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_5_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _1230_ _1575_ _1696_ _1301_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_79_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3308__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ mod.registers.r15\[6\] _3043_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _1758_ _3000_ _3001_ _2977_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6258__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4419__I _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3244__A1 mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4154__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6194__B1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3547__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__A1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3483__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3483__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6421__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ mod.registers.r15\[13\] _0810_ _0811_ mod.registers.r3\[13\] _0999_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__S _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ mod.registers.r11\[6\] _2550_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3786__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4983__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6690_ _0323_ net40 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _2507_ _2504_ _2508_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3538__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5572_ _2360_ _2458_ _2460_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1222_ _1137_ _1545_ _1319_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3408__I _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4454_ _1408_ _1476_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4948__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3405_ _0421_ _0426_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _1408_ _1409_ _1411_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6124_ mod.des.des_dout\[8\] _2848_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout81_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3336_ _3175_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6488__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _2794_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3267_ mod.funct3\[2\] _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5006_ _0911_ _1106_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5463__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5908_ _2080_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4974__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6888_ _0115_ net198 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _2350_ _2631_ _2634_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3529__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3318__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__S0 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3701__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4149__I mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5390__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5142__A1 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5443__I _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6630__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4170_ _1193_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6780__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _0038_ net157 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6742_ _0372_ net149 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3759__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ mod.registers.r14\[13\] _0980_ _0981_ mod.registers.r15\[13\] _0982_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ _0306_ net59 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3885_ mod.registers.r6\[10\] _0800_ _0792_ mod.registers.r2\[10\] _0913_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5624_ _2493_ _2494_ _2496_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6173__A3 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5381__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4184__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ mod.registers.r8\[2\] _2447_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4506_ _1151_ _1217_ _1313_ _1493_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _2365_ _2402_ _2405_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5133__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _1192_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5353__I _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4368_ _1154_ _1159_ _1293_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3695__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3695__B2 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6107_ mod.instr\[4\] _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3319_ _3141_ _3154_ _3157_ _3158_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _1326_ _1277_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__A3 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6038_ _2788_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6484__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6184__I _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3998__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6503__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4432__I _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4175__A2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6653__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3922__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5675__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3438__B2 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3610__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3610__B2 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3670_ _0501_ _0524_ mod.registers.r14\[1\] _0694_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4166__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3374__B1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ _2299_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3374__C2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A2 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ _2174_ _2251_ _2256_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4222_ _1131_ _1132_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3677__A1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4153_ _1176_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _1108_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4477__I0 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_290 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout44_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4929__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4986_ mod.pc_2\[9\] _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6725_ _0355_ net142 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _0509_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _0289_ net107 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3868_ mod.registers.r2\[11\] _0865_ _0855_ mod.registers.r9\[11\] mod.registers.r14\[11\]
+ _0820_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5607_ _2472_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6587_ _0220_ net122 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3799_ _0497_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5538_ mod.registers.r7\[13\] _2436_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__I mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ mod.registers.r6\[3\] _2391_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3668__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5811__I _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4871__B _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__I _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput18 io_in[8] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5896__A2 _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3659__A1 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3659__B2 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3241__I mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout179_I net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6699__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ mod.pc0\[1\] _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5584__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4387__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4771_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6510_ _0143_ net95 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3722_ mod.registers.r14\[0\] _0624_ _0572_ mod.registers.r6\[0\] _0750_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6441_ _3065_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5336__A1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3653_ _0546_ _0658_ _0675_ _3106_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6372_ mod.des.des_dout\[5\] net3 _3022_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3584_ mod.registers.r12\[2\] _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5323_ mod.registers.r3\[10\] _2287_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5254_ mod.registers.r2\[0\] _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ _1197_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ mod.registers.r1\[8\] _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5631__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4136_ _1163_ _0937_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6064__A2 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4067_ mod.registers.r10\[15\] _0991_ _0824_ mod.registers.r1\[15\] _0997_ mod.registers.r4\[15\]
+ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4075__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__B2 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5575__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ mod.pc_2\[7\] _1970_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6708_ _0341_ net51 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6639_ _0272_ net110 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3889__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3889__B2 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout140 net197 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout151 net154 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout162 net164 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout173 net176 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout184 net185 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout195 net196 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6841__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A3 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3813__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3416__I1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3329__B1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__C _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3236__I mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__A2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__I _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3501__B1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5941_ _2704_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6282__I _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ mod.valid0 _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _3093_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5557__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4754_ _1781_ _1778_ _0441_ _0657_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3705_ _0730_ _0507_ _0731_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5309__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4685_ _1399_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6424_ mod.registers.r15\[12\] _3055_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3636_ mod.registers.r11\[3\] _3163_ _3180_ mod.registers.r2\[3\] _0664_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__CLK net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _3012_ _3013_ _2727_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3567_ _0544_ _0590_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5306_ _2138_ _2273_ _2279_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _0539_ _2819_ _2964_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3498_ mod.funct3\[0\] _0439_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6285__A2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5237_ mod.registers.r1\[14\] _2218_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4296__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6864__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _0596_ _2121_ _2149_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4119_ _0598_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5099_ _2106_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4599__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5796__A1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3559__B1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5964__C _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4220__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4523__A2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6276__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__B2 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5446__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout211_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3970__B1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _1488_ _1496_ _1404_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ _3196_ _0434_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6478__S _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5711__A1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6140_ mod.des.des_dout\[12\] _2860_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3722__B1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3352_ mod.instr_2\[14\] _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _2709_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4278__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _2038_ _2028_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3630__S _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _2693_ _2694_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _2625_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5786_ _2336_ _2597_ _2601_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4737_ mod.ldr_hzd\[5\] _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3961__B1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4668_ _1683_ _1415_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3619_ mod.registers.r1\[3\] _3231_ _3219_ mod.registers.r4\[3\] _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6407_ _2350_ _3042_ _3045_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _1380_ _1324_ _1621_ _1622_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3713__B1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ _2999_ _3002_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6258__A2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ mod.pc_1\[10\] _2948_ _2949_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3604__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3244__A2 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4441__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3483__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6046__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__I _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6421__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ mod.registers.r8\[13\] _0813_ _0997_ mod.registers.r4\[13\] _0998_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4983__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ mod.registers.r9\[13\] _2505_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5571_ mod.registers.r8\[8\] _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3538__A3 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5932__A1 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4522_ _1404_ _1313_ _1538_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4453_ _1408_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A1 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3404_ mod.registers.r10\[7\] _0429_ _0431_ mod.registers.r7\[7\] _0432_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4384_ _1201_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6123_ mod.instr\[8\] _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5125__B _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3335_ _3138_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3424__I mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _2728_ _2795_ _2802_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout74_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3266_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _2004_ _2008_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4683__C _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5907_ _2667_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4974__A2 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6887_ _0114_ net198 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ mod.registers.r14\[5\] _2632_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ _2571_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4585__S1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__A3 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4165__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4414__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A1 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4193__A3 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5724__I _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5142__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4653__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ _0037_ net157 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4405__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _0371_ net149 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__A2 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3953_ _0518_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6290__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6672_ _0305_ net111 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3884_ mod.registers.r14\[10\] _0796_ _0786_ mod.registers.r5\[10\] _0912_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5623_ mod.registers.r9\[8\] _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5554_ _2337_ _2445_ _2449_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _1149_ _1150_ _1221_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5485_ mod.registers.r6\[9\] _2403_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5634__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _1080_ _1414_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6330__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _1249_ _0838_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3695__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6106_ _2837_ _2839_ _2840_ _2829_ _2831_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3318_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4298_ _1209_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__B _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _2789_ _2070_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3249_ mod.des.des_counter\[2\] _3095_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3383__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5544__I _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5124__A2 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3438__A2 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3610__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout124_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__B1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3374__B2 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5454__I _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ mod.registers.r2\[7\] _2252_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4221_ _0803_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6486__S _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4152_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4083_ _1110_ _1104_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4477__I1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_280 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_291 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5051__A1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _2002_ _1990_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6724_ _0354_ net144 mod.pc0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3936_ mod.registers.r7\[13\] _0962_ _0963_ mod.registers.r3\[13\] _0964_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3601__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _0288_ net105 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3867_ _0891_ _0892_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5606_ _2144_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6586_ _0219_ net130 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3798_ _0818_ _0822_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3365__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5537_ _2374_ _2435_ _2437_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5364__I _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _2340_ _2389_ _2394_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4419_ _1144_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5399_ _2340_ _2332_ _2341_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3668__A2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4708__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5290__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 io_in[9] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4002__C1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5345__A2 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__CLK net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3659__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3292__B1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A1 _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4770_ _1797_ _1794_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3595__B2 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ mod.registers.r8\[0\] _0581_ _0578_ mod.registers.r10\[0\] _0749_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ mod.des.des_dout\[16\] net19 _3061_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3652_ _0676_ _0677_ _0678_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6371_ _3023_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5184__I _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3583_ mod.registers.r8\[2\] _0490_ _0548_ mod.registers.r11\[2\] _0611_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5322_ _2194_ _2286_ _2289_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4204_ _1037_ _1058_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5184_ _2117_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _0922_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4066_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4075__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6643__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5024__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ mod.pc_2\[7\] _1970_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3586__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ _0340_ net40 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6793__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4783__B1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _0943_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4899_ _1918_ _1919_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6638_ _0271_ net110 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4212__B _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5094__I _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _0202_ net122 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3889__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4838__A1 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout130 net132 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout141 net143 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout152 net153 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout163 net164 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout174 net176 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout185 net190 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout196 net197 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3813__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4173__I _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3517__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A3 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6049__B _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3501__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3501__B2 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout191_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6666__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3252__I _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5871_ _1890_ _1828_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4822_ _0738_ _0746_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5557__A2 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4753_ mod.ldr_hzd\[8\] _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5907__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4811__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3704_ _0720_ _0721_ _0722_ _0723_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5309__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ _1708_ _1348_ _1671_ _1706_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6423_ _3036_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3635_ mod.registers.r14\[3\] _3183_ _3172_ mod.registers.r6\[3\] _0663_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3427__I _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6354_ _2997_ _2983_ _3008_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ _0593_ _0543_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5305_ mod.registers.r3\[3\] _2275_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6285_ mod.ri_3 _2820_ _2955_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3497_ _0523_ _0524_ _0443_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5236_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4296__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4258__I _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _2123_ _1967_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _1145_ _0777_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5098_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4048__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input17_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__I _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4049_ _1059_ _1071_ _1073_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__B2 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4721__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5980__C _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5720__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6689__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5484__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4039__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5787__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3970__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3970__B2 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3247__I _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _0436_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout204_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3722__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3722__B2 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5462__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _1982_ _2811_ _2813_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3282_ mod.instr_2\[10\] _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4278__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5475__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input9_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ mod.pc_2\[10\] _1106_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3486__B1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4806__I _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5923_ _2683_ mod.pc0\[9\] _2684_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4450__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ _2623_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _1828_ _1832_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5785_ mod.registers.r13\[1\] _2599_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _1761_ _3184_ _1762_ _1763_ mod.ldr_hzd\[8\] _0634_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5950__A2 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3961__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4667_ _1302_ _1296_ _1692_ _1693_ _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6406_ mod.registers.r15\[5\] _3043_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3618_ mod.registers.r7\[3\] _0431_ _3224_ mod.registers.r3\[3\] _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A2 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4505__A3 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__B _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _1139_ _1623_ _1624_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_1_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3713__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3713__B2 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6337_ _1781_ _3000_ _3001_ _1812_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3549_ mod.registers.r9\[4\] _3152_ _0576_ mod.registers.r13\[4\] _0577_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6268_ _2952_ _2947_ _2953_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5466__A1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5219_ mod.des.des_dout\[33\] _2187_ _2213_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6199_ _2896_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6378__I _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5457__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4626__I _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3530__I _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout154_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6854__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2446_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5932__A2 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4521_ _1540_ _1542_ _1548_ _1181_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _1478_ _1479_ _1339_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5696__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _1326_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6122_ _2850_ _2851_ _2852_ _2843_ _2844_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _3174_ _3155_ _3184_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ mod.pc_1\[3\] _2797_ _2799_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ mod.funct3\[1\] _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4964__C _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ _2021_ _1705_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_fanout67_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5906_ _2675_ _1926_ _1930_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_22_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _0113_ net204 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5837_ _2345_ _2631_ _2633_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5768_ _2569_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ mod.ldr_hzd\[14\] _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _2477_ _2542_ _2546_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5687__A1 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3615__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5439__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A2 _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6727__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4414__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6877__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__B1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6478__I0 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A1 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _0370_ net149 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _0624_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _0304_ net111 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3883_ mod.pc_2\[10\] _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5187__I _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4091__I _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4169__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _2474_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3916__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5553_ mod.registers.r8\[1\] _2447_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1528_ _1529_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5484_ _2360_ _2402_ _2404_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A1 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _1110_ _1414_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4366_ _1295_ _1393_ _1121_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6105_ mod.des.des_dout\[3\] _2835_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4892__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3317_ _3162_ _3142_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__I _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _1323_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4694__C _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2068_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3248_ _3095_ _3102_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__B1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A2 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _0096_ net79 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5097__I _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5825__I _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3345__I _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4332__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4885__B mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__I _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__A1 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5832__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__I _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6391__I _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4904__I _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4938__A3 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3374__A2 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__B2 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ _1163_ _1245_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _1177_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6076__A1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4477__I2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_270 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__B1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_281 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_292 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _0833_ _1987_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5051__A2 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6723_ _0353_ net148 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3935_ _3171_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _0287_ net107 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3866_ mod.registers.r12\[11\] _0893_ _0547_ mod.registers.r10\[11\] _0894_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6000__A1 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ _2481_ _2473_ _2482_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6585_ _0218_ net130 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3797_ mod.registers.r2\[8\] _0823_ _0824_ mod.registers.r1\[8\] _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5645__I _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4562__A1 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ mod.registers.r7\[12\] _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3365__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ mod.registers.r6\[2\] _2391_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4418_ _1428_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5398_ mod.registers.r5\[2\] _2334_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3522__C1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4349_ _1242_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4617__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6019_ _2774_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A3 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__B1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__C _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__C2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4069__B1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5805__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3292__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3292__B2 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5033__A2 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3720_ _3108_ _0525_ _0454_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3595__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6595__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3651_ _0667_ _0668_ _0669_ _0671_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6370_ mod.des.des_dout\[4\] net2 _3022_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3582_ mod.registers.r9\[2\] _0488_ _0493_ mod.registers.r10\[2\] _0610_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_127_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5321_ mod.registers.r3\[9\] _2287_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6297__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5252_ _2242_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4847__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ _1196_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4809__I _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4134_ _1154_ _1159_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _1082_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4967_ _1004_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6706_ _0339_ net39 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3918_ _0910_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4783__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4783__B2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4898_ _1902_ _1920_ _1903_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6637_ _0270_ net110 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3849_ _0874_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4535__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _0201_ net46 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5519_ _2351_ _2423_ _2426_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _0132_ net44 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout120 net124 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout142 net143 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout153 net154 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3510__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout164 net179 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout175 net176 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout186 net188 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout197 mod.clk net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__A2 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3577__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3329__A2 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3501__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout184_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5254__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__A3 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _2652_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5006__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4752_ _1767_ _1777_ _1778_ _1769_ _1779_ _1768_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ _0708_ _0709_ _0718_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _3121_ _1707_ _1709_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6422_ _3034_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ mod.registers.r8\[3\] _3150_ _3159_ mod.registers.r10\[3\] _0662_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _1747_ _3006_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3565_ _0591_ _0455_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5304_ _2133_ _2273_ _2278_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout97_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6284_ _2961_ _2963_ _2895_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3496_ _3229_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ mod.des.des_dout\[35\] _2159_ _2227_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__6610__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _2140_ _2167_ _2168_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ _0593_ _0543_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _1724_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5245__A2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4048_ _1059_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4274__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _2754_ _2757_ _2739_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3559__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5038__C _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3970__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6633__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3722__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3350_ mod.instr_2\[15\] _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _1879_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5475__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6783__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3486__A1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3486__B2 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A1 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3238__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _2689_ _2013_ _2016_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ _2370_ _2637_ _2642_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _1829_ _1830_ mod.valid0 _1831_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4738__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5784_ _2328_ _2597_ _2600_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ mod.ldr_hzd\[10\] _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3410__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5950__A3 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4666_ _1290_ _1305_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3961__A2 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _2345_ _3042_ _3044_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3617_ _3198_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5163__A1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _1140_ _1318_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3713__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ _2086_ _2908_ _2965_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3548_ _3139_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6267_ mod.pc_1\[9\] _2948_ _2949_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _3126_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _2113_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3477__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6198_ _2908_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5149_ _2111_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6415__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4441__A3 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6656__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4179__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6406__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6009__I1 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3640__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout147_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4196__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _1185_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _1238_ _0760_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ _3201_ _3217_ _3221_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5696__A2 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4382_ _1356_ _1357_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6121_ mod.des.des_dout\[7\] _2848_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ mod.registers.r14\[7\] _3183_ _3185_ mod.registers.r15\[7\] _3186_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _1888_ _2795_ _2801_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ _3109_ _3116_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _1731_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A1 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5905_ _2680_ _2681_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ _0112_ net204 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ mod.registers.r14\[4\] _2632_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _2501_ _2583_ _2588_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4718_ mod.ldr_hzd\[13\] _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5698_ mod.registers.r11\[1\] _2544_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4649_ _1080_ _1616_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5383__I _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5687__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ _2973_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4498__I0 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3622__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__B2 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5127__A1 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3806__I _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5678__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3689__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4102__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3541__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6821__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ mod.registers.r9\[13\] _0977_ _0978_ mod.registers.r12\[13\] _0979_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _0303_ net111 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3882_ _0906_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4305__C _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _2472_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5366__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4169__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _2329_ _2445_ _2448_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _1185_ _1359_ _1457_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4321__B _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ mod.registers.r6\[8\] _2403_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ _1408_ _1461_ _1257_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4341__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4365_ _0877_ _1292_ _1294_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6104_ _2838_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6469__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3316_ _3145_ _3153_ _3161_ _3168_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1323_ _1271_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6094__A2 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2771_ _2775_ _2779_ _2785_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3247_ _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3852__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__B2 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _0095_ net46 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ mod.registers.r13\[15\] _2617_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6799_ _0026_ net132 mod.instr_2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__A2 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4406__B _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5520__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _0437_ _0569_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6076__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _1085_ _1086_ _1087_ _1091_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_56_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4087__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__I3 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_260 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_271 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_282 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_293 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5587__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _0833_ _1987_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6722_ _0352_ net144 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3934_ _0467_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5339__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6387__I0 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3865_ _0475_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6653_ _0286_ net107 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6000__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ mod.registers.r9\[3\] _2475_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4011__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _0217_ net65 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3796_ _0483_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__B _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4562__A2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5535_ _2417_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3365__A3 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3446__I _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3770__B1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5466_ _2337_ _2389_ _2393_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4417_ _0594_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5511__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5661__I _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3522__B1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4348_ _1010_ _1218_ _1314_ _1350_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3522__C2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _1297_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4078__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _2767_ _2766_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__B1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4002__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3761__B1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4305__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A2 _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4069__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3292__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3650_ _0662_ _0663_ _0664_ _0665_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5741__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3581_ mod.registers.r5\[2\] _0423_ _3226_ mod.registers.r2\[2\] _0491_ mod.registers.r6\[2\]
+ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5320_ _2184_ _2286_ _2288_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6297__A2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4202_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ mod.des.des_dout\[29\] _2141_ _2180_ _2182_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4097__I _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _0877_ _0910_ _0947_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_96_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _1085_ _1086_ _1087_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_68_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__I _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout42_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ _1873_ _1517_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6705_ _0338_ net53 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3917_ _0605_ _0778_ _0840_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3586__A3 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4783__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ mod.pc_2\[3\] _1901_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3991__B1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6636_ _0269_ net127 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3848_ _0875_ _0868_ _0872_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6567_ _0200_ net47 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3779_ mod.registers.r9\[8\] _0805_ _0806_ mod.registers.r4\[8\] _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ mod.registers.r7\[5\] _2424_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _0131_ net44 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6288__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _2379_ _2375_ _2380_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4299__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3904__I _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout110 net111 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout121 net124 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout132 net136 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout143 net146 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout154 net155 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout165 net166 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout176 net177 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout187 net189 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout198 net199 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5799__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4471__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4471__B2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout177_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4462__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _3097_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5962__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _0501_ _0524_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4380__I _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ mod.pc_2\[1\] _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4682_ _1468_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6421_ _2370_ _3048_ _3053_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3633_ _3126_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3564_ _0513_ _0520_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6352_ _3010_ _3011_ _2727_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ mod.registers.r3\[2\] _2275_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6283_ _2092_ _1774_ _3123_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3495_ mod.instr_2\[3\] _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _2190_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5165_ mod.registers.r1\[6\] _2146_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4116_ _1138_ _1141_ _1143_ _1139_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_68_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6256__B _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4047_ _1074_ _0986_ _1070_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5953__A1 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _1036_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ _0252_ net125 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4508__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6585__CLK net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4444__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__B _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4747__A2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3544__I _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A1 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3280_ mod.instr_2\[11\] _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3486__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _2669_ _1995_ _2692_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ mod.registers.r14\[11\] _2638_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6188__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6188__B2 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ net13 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A1 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ mod.registers.r13\[0\] _2599_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4734_ _1750_ _3136_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3410__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _0947_ _1167_ _1304_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6404_ mod.registers.r15\[4\] _3043_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3616_ _0621_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5163__A2 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _1608_ _1225_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6335_ _2973_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3547_ mod.registers.r14\[4\] _0469_ _3164_ mod.registers.r11\[4\] _0575_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _2005_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3478_ mod.pc_2\[5\] _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5217_ _1970_ _2190_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6197_ _1804_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _2087_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6415__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5079_ mod.rd_3\[3\] _2083_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__I _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5844__I _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5154__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4195__I _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4417__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__A2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__B _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6600__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4450_ _1368_ _0769_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6750__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3401_ _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4381_ _1165_ _0954_ _0922_ _1045_ _1338_ _1207_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_6120_ _2663_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3332_ _3184_ _3138_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6051_ mod.pc_1\[2\] _2797_ _2799_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3263_ _3112_ _3115_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _2019_ _1887_ _2001_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3864__C1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4833__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _2678_ mod.pc0\[3\] _0003_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6884_ _0111_ net202 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3631__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5835_ _2625_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3449__I _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5766_ mod.registers.r12\[11\] _2584_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4717_ mod.ldr_hzd\[12\] _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5697_ _2470_ _2542_ _2545_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4648_ _1616_ _0985_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _1593_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6318_ _2985_ _2987_ _2981_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6249_ _2892_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4647__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4498__I1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3622__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6773__CLK net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4430__S0 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4102__A3 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3861__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5749__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _0516_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _0908_ _0901_ _0904_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3269__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _2183_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4169__A3 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5551_ mod.registers.r8\[0\] _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _1210_ _1453_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6315__A1 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _2390_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _1165_ _1155_ _1249_ _1460_ _1269_ _1266_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4877__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4364_ _1349_ _1354_ _1385_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6103_ _2662_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4828__I _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3315_ mod.registers.r11\[7\] _3164_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _1242_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4629__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3246_ _3100_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout72_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _2714_ _2786_ _2787_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4049__B _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6646__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6796__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6867_ _0094_ net75 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5818_ _2381_ _2616_ _2620_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5357__A2 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6798_ _0025_ net165 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5749_ _2571_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6306__A1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A1 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3828__C1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5569__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A2 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3359__A1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6519__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4859__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__B _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6669__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4080_ _1094_ _1105_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A1 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4584__S _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_250 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_261 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_272 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_283 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_294 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5036__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _1843_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6721_ _0351_ net143 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3933_ mod.registers.r13\[13\] _0959_ _0960_ mod.registers.r6\[13\] _0961_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6652_ _0285_ net121 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6387__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ mod.registers.r5\[11\] _0559_ _0806_ mod.registers.r4\[11\] _0858_ mod.registers.r8\[11\]
+ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5603_ _2137_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _0216_ net65 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3795_ _0477_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__I _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _2415_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3770__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3770__B2 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5465_ mod.registers.r6\[1\] _2391_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4416_ _1442_ _1443_ _1145_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5511__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _2132_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3522__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3522__B2 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4347_ _1367_ _1331_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3462__I _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _1163_ _0937_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5275__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ mod.pc\[10\] _2030_ _1890_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4507__B _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5389__I _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6224__B1 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3589__B2 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4002__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3761__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3761__B2 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__B1 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4931__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout122_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _0606_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6491__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4201_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5181_ _2152_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _0832_ _0839_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5257__A1 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4063_ _1088_ _1089_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4965_ _1728_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__I mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4841__I _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6704_ _0337_ net106 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3916_ _0877_ _0910_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3440__B1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ mod.pc_2\[3\] _1901_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6635_ _0268_ net127 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3991__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3847_ _0841_ _0853_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3991__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6834__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5193__B1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _0199_ net47 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5732__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3778_ _3218_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5517_ _2346_ _2423_ _2425_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6497_ _0130_ net43 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5672__I _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5448_ mod.registers.r5\[13\] _2376_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4299__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout100 net101 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout111 net112 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5379_ mod.registers.r4\[14\] _2323_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout122 net124 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout133 net134 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout144 net145 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout155 net156 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout166 net169 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5248__A1 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout177 net178 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout188 net189 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4471__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3431__B1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3982__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5723__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3734__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A3 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3830__I _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6707__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6857__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0613_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3701_ _3199_ _0689_ _0702_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4681_ _3121_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6420_ mod.registers.r15\[11\] _3049_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3632_ _0645_ _0648_ _0656_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3725__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ _2997_ _2977_ _3008_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5492__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3563_ mod.pc_2\[5\] _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ _2127_ _2273_ _2277_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6282_ _2804_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3494_ _0499_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5478__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _2006_ _2163_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3489__B1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4150__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ _1142_ _1140_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _2087_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _3194_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _2721_ _2729_ _2747_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4948_ _0411_ _0433_ _1915_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4879_ _1902_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6618_ _0251_ net125 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3716__A1 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3716__B2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6549_ _0182_ net72 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4516__I0 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__B1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3891__B1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4435__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ _2668_ mod.pc0\[8\] _2673_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3643__B1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5851_ _2367_ _2637_ _2641_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6188__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4199__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ mod.valid2 _1827_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5782_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5935__A2 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ mod.ldr_hzd\[11\] _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4664_ _1291_ _0942_ _0949_ _1295_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5699__A1 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _3036_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3615_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4595_ _1221_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3735__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6334_ _2651_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3546_ mod.registers.r15\[4\] _0518_ _0509_ mod.registers.r1\[4\] _0574_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _0779_ _2947_ _2951_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ _0473_ _0498_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_88_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4123__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _2062_ _2121_ _2196_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6196_ _2889_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4674__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5871__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5147_ _0591_ _2121_ _2149_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5078_ _2081_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _1053_ _1054_ _1055_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3634__B1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__I _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5926__A2 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6552__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4665__A2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4476__I _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__C _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4417__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3555__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout202_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ _0412_ _0414_ _0427_ _3205_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4380_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4353__B2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ _3162_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _2720_ _2795_ _2800_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3262_ _3114_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ mod.pc\[10\] _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__C2 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5605__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4408__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A2 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _2675_ _1908_ _1912_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_53_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6883_ _0110_ net204 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _2623_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6030__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _2499_ _2583_ _2587_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4716_ net14 _1741_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5696_ mod.registers.r11\[0\] _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _1121_ _1171_ _1674_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3465__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4344__A1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4578_ _1469_ _1599_ _1600_ _1601_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_1_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6317_ _2970_ _2986_ _2979_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3529_ mod.registers.r6\[4\] _0491_ _0484_ mod.registers.r4\[4\] _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _2657_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3414__B _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _2891_ _2894_ _2895_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__I _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4032__B1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4583__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3630__I0 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6324__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4335__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4430__S1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A3 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__A2 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout152_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _0883_ _0888_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6598__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4574__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _1243_ _1409_ _1256_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5481_ _2388_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4432_ _0473_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4877__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4363_ _1388_ _1389_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6102_ mod.instr\[3\] _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3314_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _1229_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5826__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ mod.pc\[12\] _2714_ _2751_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3245_ _3099_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _0093_ net75 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6003__A1 _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ mod.registers.r13\[14\] _2617_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _0024_ net165 mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5748_ _2569_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ mod.registers.r10\[11\] _2529_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6306__A2 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4868__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__I _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5817__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3828__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A2 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A2 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__A1 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6740__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5808__A1 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4087__A3 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_240 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_251 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_262 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_273 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_284 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_295 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5036__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _0861_ _0867_ _1853_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6720_ _0350_ net142 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ _0572_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4795__A1 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6651_ _0284_ net121 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3863_ mod.registers.r15\[11\] _0558_ _0551_ mod.registers.r7\[11\] _0859_ mod.registers.r3\[11\]
+ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4613__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5602_ _2479_ _2473_ _2480_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4547__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ _0215_ net63 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3794_ mod.registers.r5\[8\] _0819_ _0821_ mod.registers.r14\[8\] _0822_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5533_ _2371_ _2429_ _2434_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3770__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5464_ _2329_ _2389_ _2392_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3507__C1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4415_ _1200_ _1273_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5395_ _2337_ _2332_ _2338_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4346_ _1370_ _1372_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3522__A2 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _1167_ _1304_ _0947_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6016_ _2771_ _2768_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3825__A3 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6224__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6224__B2 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3589__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _0076_ net208 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3761__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__I _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5266__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5018__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__B2 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6636__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout115_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ _1184_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4701__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _1901_ _2153_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6786__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4131_ _1156_ _1157_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5257__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4062_ mod.registers.r8\[15\] _0971_ _0981_ mod.registers.r15\[15\] _1090_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ mod.pc0\[8\] _1835_ _1983_ _1857_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6703_ _0336_ net103 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3915_ _0938_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4895_ _0871_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3440__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3440__B2 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6634_ _0267_ net127 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3846_ _0854_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3991__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6565_ _0198_ net45 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3777_ _0488_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5516_ mod.registers.r7\[4\] _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6496_ _0129_ net99 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5447_ _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3473__I _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5378_ _2225_ _2322_ _2325_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout101 net114 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout134 net135 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4329_ _1232_ _1240_ _1269_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout145 net146 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout156 net196 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout167 net169 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5248__A2 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout178 net179 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout189 net190 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4456__B1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6509__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3431__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3648__I mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3431__B2 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3734__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3498__A1 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5239__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4428__B _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3670__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3558__I _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _0539_ _0502_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _1288_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _0538_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6350_ _1746_ _3006_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3562_ _0567_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3725__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4610__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5301_ mod.registers.r3\[1\] _2275_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ net20 _2959_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3493_ _0506_ _0507_ _0513_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5478__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _2107_ _2073_ _2163_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3489__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3489__B2 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ mod.des.des_dout\[27\] _2159_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6427__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ _0619_ _0620_ _0642_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5094_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4438__B1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6109__I _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4045_ _0441_ _1072_ _3165_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1960_ _1962_ _1977_ _1978_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5402__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4947_ _1967_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _0766_ _1880_ _1735_ _1863_ _1881_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6617_ _0250_ net131 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5166__A1 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ mod.registers.r15\[9\] _0558_ _0555_ mod.registers.r12\[9\] _0551_ mod.registers.r7\[9\]
+ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4913__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _0181_ net63 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6479_ _3087_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5469__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4516__I1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3931__I _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4248__B _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5641__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3652__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3652__B2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__A1 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__I0 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3378__I _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3404__B2 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3891__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout182_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5768__I _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3643__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3643__B2 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ mod.registers.r14\[10\] _2638_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4801_ _1725_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4199__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _2595_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4732_ _1758_ _1759_ _3155_ _0711_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4663_ _3132_ _1673_ _1675_ _1682_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3614_ _0622_ _0522_ _0630_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6402_ _3034_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4594_ _1608_ _1620_ _1389_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6333_ _2996_ _2998_ _2993_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3545_ mod.registers.r4\[4\] _0570_ _0571_ mod.registers.r2\[4\] _0572_ mod.registers.r6\[4\]
+ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ mod.pc_1\[8\] _2948_ _2949_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3476_ _0500_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _2123_ _2047_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5320__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _2899_ _2906_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5146_ _2129_ _1933_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5077_ _1809_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4028_ mod.registers.r3\[14\] _0963_ _0972_ mod.registers.r2\[14\] _1056_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3634__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3634__B2 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _2650_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3398__B1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5139__A1 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4531__B _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__I _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5311__A1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5378__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4889__B1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _3178_ _3179_ _3138_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__A1 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3261_ _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ mod.pc0\[10\] _1889_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_112_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__B2 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3616__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _2676_ _2679_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6882_ _0109_ net212 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5369__A1 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _2342_ _2624_ _2630_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6030__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ mod.registers.r12\[10\] _2584_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ net15 _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5695_ _2543_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4646_ _1078_ _1128_ _1170_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_163_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5541__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4577_ _1441_ _1314_ _1483_ _1603_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6316_ _1799_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ mod.registers.r8\[4\] _0490_ _0555_ mod.registers.r12\[4\] _0556_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _0622_ _2658_ _2939_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3459_ _0422_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3481__I _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3414__C mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6178_ _2659_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _2108_ _1896_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5072__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4032__B2 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3630__I1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4335__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5532__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3689__A4 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5599__A1 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout145_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4023__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__B2 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3377__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4500_ _1205_ _1526_ _1527_ _1407_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5480_ _2357_ _2396_ _2401_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4431_ _1377_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5523__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4362_ _1386_ _1387_ _1350_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6101_ _2834_ _2664_ _2836_ _2829_ _2831_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3313_ mod.instr_2\[1\] _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4293_ _1316_ _1319_ _1320_ _0906_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3244_ mod.des.des_counter\[0\] mod.des.des_counter\[1\] _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _2783_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6542__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6865_ _0092_ net56 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__I mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _2378_ _2616_ _2619_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4014__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6796_ _0023_ net166 mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5747_ _2481_ _2570_ _2576_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4565__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6692__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3773__B1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _2499_ _2528_ _2532_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4317__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0505_ _1655_ _1654_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3828__B2 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__I _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4005__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__B1 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3819__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_230 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4492__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_241 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_252 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6565__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_263 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_274 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_285 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_296 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5036__A3 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4980_ _1873_ _1427_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3931_ _0576_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4795__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3497__S _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _0283_ net123 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _0878_ _0780_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ mod.registers.r9\[2\] _2475_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4547__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _0214_ net63 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3793_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3755__B1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5532_ mod.registers.r7\[11\] _2430_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5463_ mod.registers.r6\[0\] _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3507__B1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4414_ _1432_ _1437_ _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5394_ mod.registers.r5\[1\] _2334_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _1189_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4276_ _1154_ _1159_ _1303_ _1293_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6015_ _2756_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3286__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4076__B _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6291__B _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _0075_ net205 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _0409_ net166 mod.instr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3934__I _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4710__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__CLK net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4765__I mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3277__A2 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4226__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__B1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6220__I _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4701__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4130_ _1155_ _0450_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ mod.registers.r4\[15\] _0974_ _0972_ mod.registers.r2\[15\] _0975_ mod.registers.r11\[15\]
+ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _1982_ _1889_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _0335_ net105 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3914_ _0941_ _0931_ _0936_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4894_ mod.pc_2\[4\] _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3440__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _0266_ net125 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5717__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3845_ _0868_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6564_ _0197_ net56 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3776_ _0645_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5515_ _2417_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3754__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6495_ _0128_ net100 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5446_ _2224_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6730__CLK net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ mod.registers.r4\[13\] _2323_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout102 net104 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3900__B1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout124 net129 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout135 net136 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4328_ _1355_ _1197_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout146 net156 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout157 net196 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout168 net169 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout179 net195 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4259_ _1114_ _1115_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6880__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__B2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3929__I mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6305__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3431__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5708__A1 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A3 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4695__A1 _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4709__B _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__A3 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4447__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3670__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__I _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3630_ mod.funct7\[0\] _0657_ _0442_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6753__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3561_ _0568_ _0569_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3725__A3 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _2116_ _2273_ _2276_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6280_ _2959_ _2960_ _2895_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3492_ _0514_ _0515_ _0517_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5231_ _2211_ _2225_ _2226_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4686__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3489__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _2159_ _2161_ _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ _0770_ _0771_ _1139_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5093_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _3106_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4989__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3661__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout40_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5938__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _2748_ _2749_ _1977_ _1978_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6125__I _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1731_ _1670_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4610__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4877_ _0766_ _1880_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6616_ _0249_ net41 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ mod.registers.r5\[9\] _0559_ _0806_ mod.registers.r4\[9\] _0855_ mod.registers.r9\[9\]
+ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5166__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6547_ _0180_ net48 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3716__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3759_ mod.registers.r5\[8\] _0786_ _0677_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4913__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6478_ mod.des.des_dout\[32\] net4 _3084_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _2364_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6418__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6626__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3652__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4601__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4452__I1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3404__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3340__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3891__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4515__S1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout175_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3643__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _2596_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _3178_ _1749_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _1286_ _1079_ _1672_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4621__C _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _2342_ _3035_ _3041_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3613_ _0631_ _0633_ _0638_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4593_ _1608_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6332_ _2997_ _2986_ _2978_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3544_ _3172_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4108__B1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _0596_ _2947_ _2950_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3475_ _0502_ mod.funct3\[1\] _0445_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4659__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ _2102_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6194_ _1793_ _2900_ _2904_ mod.instr\[4\] _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_fanout88_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _0440_ _2082_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5084__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__I _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ mod.registers.r8\[14\] _0971_ _0968_ mod.registers.r10\[14\] _1055_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3634__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _2737_ _2738_ _2739_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3398__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__B2 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _1452_ _1485_ _1858_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4812__B mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6336__A1 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4103__I _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3570__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4114__A3 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4259__B _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__I _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4822__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3610__C _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3389__A1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5109__I _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4889__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__S0 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4889__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3561__A1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3260_ mod.instr_2\[0\] _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3313__A1 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__D _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3616__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _2678_ mod.pc0\[2\] _0003_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3299__I _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6881_ _0108_ net202 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5832_ mod.registers.r14\[3\] _2626_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4577__B1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _2497_ _2583_ _2586_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4632__B _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4714_ mod.ins_ldr_3 mod.valid_out3 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6403__I _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _2540_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ _1079_ _1302_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4576_ _1440_ _1318_ _1221_ _0776_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6315_ _1756_ _2974_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _3210_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6246_ mod.pc_1\[2\] _2936_ _2822_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3458_ _0476_ _0479_ _0482_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_103_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _2092_ _2893_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3389_ _3201_ _3216_ _3211_ _3220_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5128_ _2103_ _2133_ _2134_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _2059_ _1691_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_73_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A1 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4032__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__I _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6814__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5532__A2 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5048__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4559__B1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4023__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout138_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6494__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _0954_ _1163_ _0985_ _1045_ _1368_ _1355_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _1124_ _3130_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6100_ mod.des.des_dout\[2\] _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3312_ _3110_ _3113_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4292_ _1222_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5287__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _2054_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3243_ _3098_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6864_ _0091_ net89 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ mod.registers.r13\[13\] _2617_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6795_ _0022_ net165 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6837__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ mod.registers.r12\[3\] _2572_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5762__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3773__A1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3773__B2 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ mod.registers.r10\[10\] _2529_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4628_ _1654_ _0505_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4559_ _1285_ _1583_ _1584_ _1380_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__A1 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ _0693_ _2924_ _2927_ mod.instr\[16\] _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3828__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3461__B1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4005__A2 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6043__I _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__B1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5882__I _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_220 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4447__B _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_231 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_242 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__B1 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_253 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_264 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_275 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_286 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_297 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3930_ _0780_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4795__A3 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ _0883_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ _2132_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6580_ _0213_ net51 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3792_ _3213_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5744__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3755__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5531_ _2368_ _2429_ _2433_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3755__B2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5792__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5462_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3507__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4413_ _1438_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3507__B2 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5393_ _2336_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4201__I _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4344_ _1371_ _1262_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4275_ _0948_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout70_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6014_ mod.pc\[10\] _2763_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5680__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3286__A3 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6128__I mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5032__I _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__C _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _0074_ net205 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _0408_ net166 mod.instr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3746__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5729_ _2507_ _2561_ _2564_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5499__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__I _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__I _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__B _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4781__I mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3985__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__B2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3397__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5726__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ mod.registers.r13\[15\] _0959_ _0980_ mod.registers.r14\[15\] _1088_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6682__CLK net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ mod.pc\[8\] _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3913_ mod.pc_2\[10\] _3127_ _0939_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3976__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6701_ _0334_ net106 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4893_ _3094_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6632_ _0265_ net82 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3844_ _0763_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5717__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3728__A1 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _0196_ net57 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3728__B2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3775_ _0779_ _0780_ _0790_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_164_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5514_ _2415_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _0127_ net98 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5445_ _2374_ _2375_ _2377_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5376_ _2217_ _2322_ _2324_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout103 net104 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4866__I _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3900__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3361__C1 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _1338_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout114 net139 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout125 net128 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3900__B2 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout136 net137 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout147 net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout158 net159 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout169 net178 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5653__A1 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _1215_ _1216_ _1179_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3664__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3719__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4550__B _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6555__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A1 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__I mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5644__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4998__A3 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3670__A3 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5400__I _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4016__I mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout120_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6231__I _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ _0573_ _0580_ _0584_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_6_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ mod.registers.r14\[5\] _0469_ _0518_ mod.registers.r15\[5\] _0519_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5230_ mod.registers.r1\[13\] _2218_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5161_ _0503_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__B1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ _0681_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ _2090_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4043_ _3196_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3497__I0 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ mod.pc\[7\] _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4945_ _1875_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4071__B1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4876_ _0830_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6615_ _0248_ net41 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3827_ _0424_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6141__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6546_ _0179_ net45 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3758_ _3156_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6477_ _3086_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3689_ _0714_ _3136_ mod.registers.r2\[1\] _0712_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5428_ _2193_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5874__A1 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5359_ mod.registers.r4\[6\] _2311_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3885__B1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6316__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5220__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__B _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6354__A2 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__A2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5890__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4117__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3340__A2 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6226__I _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout168_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4730_ mod.ldr_hzd\[9\] _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4661_ _1334_ _1685_ _1687_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3585__I _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ mod.registers.r15\[3\] _3037_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6870__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4356__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3612_ mod.registers.r9\[2\] _0639_ _0582_ mod.registers.r3\[2\] _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _0772_ _1138_ _0770_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _2908_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3543_ _3180_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4108__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ mod.pc_1\[7\] _2948_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4108__B2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3474_ mod.instr_2\[4\] _0501_ _0442_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5856__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _2176_ _2209_ _2210_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6193_ _2899_ _2905_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _2111_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5075_ mod.rd_3\[2\] _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3619__B1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6281__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4026_ mod.registers.r15\[14\] _0981_ _0978_ mod.registers.r12\[14\] _1054_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6136__I _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6033__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _2704_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3398__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _3102_ _1947_ _1949_ _1917_ _1950_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__3495__I mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _1879_ _1883_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4347__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _0162_ net39 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5847__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3858__B1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3873__A3 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A1 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4822__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__B1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6893__CLK net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4338__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3561__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5838__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3313__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4185__B _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6880_ _0107_ net202 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _2339_ _2624_ _2629_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A1 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ mod.registers.r12\[9\] _2584_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4577__B2 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4713_ _1072_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _2541_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4329__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _1078_ _1042_ _1048_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4575_ _1505_ _1602_ _1235_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3526_ mod.registers.r14\[4\] _0481_ _0478_ mod.registers.r3\[4\] _0554_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6314_ _2982_ _2984_ _2981_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5829__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _0707_ _2658_ _2938_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3457_ mod.registers.r1\[6\] _0483_ _0484_ mod.registers.r4\[6\] _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4501__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6176_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6766__CLK net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3388_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5127_ mod.registers.r1\[2\] _2118_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6254__A1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ _1875_ _2060_ _2061_ _1851_ _2072_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_55_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4804__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _0456_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4568__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4784__I _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5048__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4559__B2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6440__S _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout200_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1350_ _1386_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4731__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6789__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3311_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ mod.pc\[12\] _1857_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3242_ _3097_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4798__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ _0090_ net57 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5814_ _2373_ _2616_ _2618_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _0021_ net158 mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ _2479_ _2570_ _2575_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3773__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ _2497_ _2528_ _2531_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4627_ _0594_ _1444_ _1428_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4558_ _3119_ _1142_ _1585_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3509_ _0532_ _0536_ _3108_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4489_ _1487_ _1497_ _1498_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_1_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _2923_ _2928_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _2877_ _2875_ _2878_ _2879_ _2880_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6227__B2 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4789__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3997__C1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3461__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3461__B2 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__B2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3683__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4713__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5269__A2 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_221 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4447__C _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6218__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_232 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6218__B2 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_243 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4492__A3 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_254 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_265 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_276 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_287 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_298 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4795__A4 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout150_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _0884_ _0885_ _0886_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_32_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ _0487_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3755__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ mod.registers.r7\[10\] _2430_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5461_ _2387_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _0775_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3507__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _2126_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ _1204_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _2764_ _2769_ _2660_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5680__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout63_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3691__A1 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6480__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4640__B1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3768__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6144__I mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _0073_ net205 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _0407_ net168 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4243__I0 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3989_ _1013_ _1014_ _1015_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_10_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ mod.registers.r11\[13\] _2562_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5659_ mod.registers.r10\[3\] _2517_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5932__B _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6319__I _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A1 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6471__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3434__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A2 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A2 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4934__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__B1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4961_ _1966_ _1968_ _1969_ _1917_ _1981_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4473__I0 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _0333_ net127 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3912_ _0917_ _0918_ _0919_ _0920_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4892_ _0553_ _0561_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _0264_ net82 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5178__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3843_ _0869_ _0564_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4921__B mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3728__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3774_ _0793_ _0795_ _0798_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6562_ _0195_ net58 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5513_ _2343_ _2416_ _2422_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5308__I _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6493_ _0126_ net100 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ mod.registers.r5\[12\] _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4153__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5350__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ mod.registers.r4\[12\] _2323_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3361__B1 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout104 net113 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4326_ _1350_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3900__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout115 net119 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3361__C2 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout126 net128 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout137 net138 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6139__I mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout148 net155 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5102__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4257_ _3118_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout159 net164 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4188_ _3122_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3664__A1 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__B2 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5169__A1 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6829_ _0056_ net191 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4122__I _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5888__I _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3655__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3670__A4 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4907__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3490_ _3185_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4967__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3894__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ _0674_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3894__B2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5091_ _2097_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _0986_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3646__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__B1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3497__I1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ _2746_ _2706_ _2752_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4207__I _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1876_ _1951_ _1952_ _1917_ _1965_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4071__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4071__B2 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _1727_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__I _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _0247_ net44 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3826_ _0841_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _0178_ net64 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5571__A1 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3757_ mod.registers.r13\[8\] _0784_ _0586_ mod.registers.r12\[8\] _0785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3582__B1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6476_ mod.des.des_dout\[31\] net3 _3084_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3688_ _3147_ _0635_ mod.registers.r4\[1\] _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5323__A1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4126__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _2360_ _2361_ _2363_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5358_ _2157_ _2310_ _2313_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3885__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3885__B2 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5289_ _2231_ _2263_ _2267_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3637__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6522__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5562__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6672__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4117__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A1 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6000__C _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5411__I _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4660_ _1077_ _1225_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _3151_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5553__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _1412_ _1341_ _1615_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6330_ _1767_ _2988_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3542_ _3176_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4108__A2 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _2814_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3473_ _3232_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5212_ mod.registers.r1\[11\] _2185_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ mod.instr_2\[3\] _2900_ _2904_ mod.instr\[3\] _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5143_ _2140_ _2145_ _2147_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _2081_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3619__B2 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4025_ mod.registers.r9\[14\] _0977_ _0967_ mod.registers.r5\[14\] _1053_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6545__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _2730_ _2736_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_40_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _3098_ _1933_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3776__I _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6152__I _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _1862_ _1877_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6336__A3 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3809_ _0833_ _0834_ _0835_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4789_ mod.instr_2\[6\] _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6528_ _0161_ net96 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4752__C1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _3075_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4400__I _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3858__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3858__B2 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6272__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A2 _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A1 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3389__A3 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3794__B1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__B1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5406__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__S _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__A2 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout180_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5141__I _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ mod.registers.r14\[2\] _2626_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4026__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4026__B2 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5774__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5761_ _2493_ _2583_ _2585_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3596__I _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4712_ _3116_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5692_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4329__A2 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _1392_ _1631_ _1652_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5526__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ _1339_ _1512_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _2970_ _2983_ _2979_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3525_ _0549_ _0550_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6244_ mod.pc_1\[1\] _2936_ _2822_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout93_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ _3218_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _2656_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3387_ _0413_ _0414_ _3209_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6254__A2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6147__I mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _3100_ _2068_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_55_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4008_ _0524_ _1034_ _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5986__I mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4568__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ _1837_ _1839_ mod.pc\[2\] _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__B _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5517__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3528__B1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6057__I _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3464__C1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4008__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4559__A2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3767__B1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5508__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__I _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3310_ _3146_ _3148_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_99_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _3118_ _1317_ _1219_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3241_ mod.des.des_counter\[0\] _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4908__C _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__B _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4247__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _0089_ net59 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3470__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ mod.registers.r13\[12\] _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5747__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _0020_ net158 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ mod.registers.r12\[2\] _2572_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ mod.registers.r10\[9\] _2529_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ _1147_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6172__B2 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6733__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4557_ _1216_ _1142_ _0771_ _1180_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3508_ _0533_ _0534_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4488_ _1220_ _1499_ _1503_ _1504_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_103_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6227_ _0501_ _2924_ _2927_ mod.instr\[15\] _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3439_ _3187_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6883__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _2650_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5109_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6089_ mod.des.des_dout\[0\] _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__B1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3997__C2 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3461__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3964__I _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_222 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_233 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_244 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_255 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_266 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_277 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_288 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_299 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3988__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout143_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ mod.registers.r6\[8\] _0816_ _0555_ mod.registers.r12\[8\] mod.registers.r13\[8\]
+ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__6756__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5460_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6154__B2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4411_ _0589_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5901__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2329_ _2332_ _2335_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4342_ _1270_ _1274_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4273_ _1120_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4638__C _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _2765_ _2766_ _2768_ _2757_ _2713_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

