* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_79_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3140__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3155_ _2421_ _2374_ _2423_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3086_ _2383_ _2315_ _2175_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout56_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2953__I mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3988_ _2264_ _0972_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3784__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2939_ _2217_ _2226_ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4156__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ mod.des.des_dout\[25\] _1573_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__B1 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3198__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2796__I1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3370__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5183__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2720__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ mod.pc_1\[11\] _1833_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4622__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ _0921_ _0885_ _0805_ _0884_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _1651_ _1784_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3842_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3189__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3773_ _0781_ _0782_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4925__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2936__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2787__I1 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ mod.des.des_dout\[14\] net10 _2059_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2655_ _2164_ _2023_ _2019_ mod.instr\[9\] _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _0261_ net145 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2586_ _0003_ _1481_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3361__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ mod.pc\[8\] _1292_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout105 net108 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout116 net132 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout127 net130 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout138 net141 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4256_ mod.pc_2\[0\] _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3113__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3207_ mod.registers.r4\[3\] _2228_ _2224_ mod.registers.r3\[3\] _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4187_ _2253_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2711__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3138_ _2148_ _2435_ _2426_ mod.registers.r2\[1\] _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3069_ _2230_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3728__B _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2778__I1 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3019__I _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2858__I _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3104__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2702__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3689__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__C _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4110_ _0881_ _1118_ _1119_ _0920_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5090_ mod.instr\[3\] _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4041_ _0708_ _0654_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _1388_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2606__B1 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__A2 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ _1594_ mod.registers.r6\[6\] _1770_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3548__B _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3825_ _2309_ _0678_ _2527_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3756_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2707_ _2052_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3687_ _0437_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4206__S0 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2638_ _2013_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3283__B _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3334__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ _0244_ net57 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2569_ mod.instr\[15\] _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3885__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2688__A3 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _1248_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _0175_ net107 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4239_ _1204_ _2129_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2860__A3 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2789__S _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4117__A3 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3325__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5221__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5371__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5002__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3610_ _2267_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3939__I0 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _1266_ _1575_ _1578_ _1538_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3541_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2699__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3472_ _0440_ mod.registers.r3\[8\] _2223_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _0101_ net73 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5142_ _0032_ net59 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5069__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4024_ _0569_ _0843_ _0791_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3095__A3 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4292__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2961__I _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4926_ mod.ri_3 _1800_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _1660_ mod.registers.r6\[0\] _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _0814_ _0730_ _0817_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4788_ _1581_ mod.registers.r4\[5\] _1728_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3739_ _2526_ _2528_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_109_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4807__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5244__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4283__A2 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2871__I _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3794__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2597__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__S _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4594__I0 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3849__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3651__B _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4274__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2972_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3785__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _0478_ _1674_ _1680_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2588__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _1625_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3826__B _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5117__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4573_ _2523_ _1545_ _1546_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3524_ _2190_ _0516_ _0530_ _2340_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3455_ mod.registers.r1\[8\] _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3117__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout86_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3304__A4 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3386_ _2469_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5125_ _0015_ net36 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2956__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _1918_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4265__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _2263_ _0895_ _1004_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_84_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A2 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4909_ mod.rd_3\[0\] _1800_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3240__A3 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__B _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4256__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2742__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3240_ _2211_ mod.registers.r3\[7\] _2359_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3152__C1 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4495__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3171_ _2202_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4247__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3207__B1 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4940__B _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3222__A3 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2886_ _2178_ _2182_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4625_ _1582_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2981__A2 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _2444_ _1545_ _1546_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_116_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3930__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3507_ _2137_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _0427_ _0434_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ mod.funct7\[2\] _2517_ _2274_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4486__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _2149_ _2153_ _2176_ mod.registers.r2\[9\] _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ mod.instr\[8\] _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__S _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5039_ mod.pc\[10\] _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3461__A3 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4410__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput20 net20 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4477__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2596__I _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_201 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_212 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_223 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_234 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_245 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_256 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_267 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_278 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_289 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3988__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__I0 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ _1565_ _2068_ _2072_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout136_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2671_ mod.funct7\[0\] _2030_ _2010_ mod.instr\[15\] _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _1416_ _1083_ _1359_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3912__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _1250_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3223_ _2331_ _2332_ _2519_ mod.registers.r2\[3\] _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3140__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3154_ _2450_ _2451_ _2131_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5305__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3085_ _2166_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3979__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout49_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2651__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__B _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3987_ _0632_ _0989_ _0991_ _0510_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2938_ mod.registers.r4\[15\] _2229_ _2235_ mod.registers.r1\[15\] _2236_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3286__B _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _2166_ _2151_ _2143_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4156__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _1595_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4156__B2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3903__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4896__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4539_ _1532_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3040__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2642__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__B2 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__B _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3198__A2 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3370__A2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5328__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3215__I mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A2 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3425__A3 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4622__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3910_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4890_ _1645_ _1774_ _1790_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3841_ _0312_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3189__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3772_ _0552_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2936__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2723_ _2061_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4138__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2654_ _1796_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5373_ _0260_ net147 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2585_ _1985_ _1458_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _1321_ _1325_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_113_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout106 net107 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout117 net118 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4255_ _0658_ _0311_ _0295_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout139 net141 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3113__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3206_ mod.registers.r5\[3\] _2200_ _2209_ mod.registers.r2\[3\] _2215_ mod.registers.r6\[3\]
+ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_4186_ _0742_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3137_ _2151_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2872__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3068_ mod.registers.r7\[0\] _2365_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3795__I _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4129__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3352__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3104__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2874__I _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4368__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5150__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5096__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ _0795_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4485__B _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4843__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1420_ _1826_ _1821_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2606__A1 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2606__B2 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _1781_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3824_ _0828_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5020__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3755_ _0670_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2706_ mod.des.des_dout\[6\] net2 _2049_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3686_ _0690_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4206__S1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2637_ _2125_ _1797_ _1930_ mod.instr\[2\] _1809_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3334__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5356_ _0243_ net72 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2568_ _1976_ _1970_ _1977_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _2122_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _0174_ net106 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4238_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_87_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _0899_ _0908_ _0693_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4047__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5173__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3325__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__I1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3013__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ _2452_ _2454_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4761__A1 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3471_ _2231_ _0398_ _2233_ mod.registers.r4\[8\] _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5210_ _0100_ net76 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _0031_ net41 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__C _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _1507_ _1350_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ _0540_ _0919_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3095__A4 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4925_ _1240_ _1799_ _1814_ _1815_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4856_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _0733_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4787_ _1718_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3555__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3738_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3669_ _0677_ _0679_ _2449_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3307__A2 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4504__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _0226_ net148 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4409__I _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2818__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3243__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3794__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4594__I1 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A3 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3932__B _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3651__C _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4482__C _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2971_ _2191_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3234__A1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _1609_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3785__A2 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4641_ _1624_ mod.registers.r1\[10\] _1554_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4734__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _1556_ _1391_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3523_ _0518_ _0530_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4003__B _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3454_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4498__B1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3385_ mod.registers.r7\[9\] _2219_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5124_ _0014_ net40 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout79_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5055_ _0003_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ _0900_ _0853_ _1014_ _0694_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3473__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2972__I _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4899__I _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4839_ _0467_ _1754_ _1760_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3528__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__B _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5211__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3700__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3464__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A1 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4716__A1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3152__B1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3152__C2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ mod.registers.r2\[2\] _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2750__I0 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3470__A4 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4255__I0 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3207__B2 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2954_ _2251_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3222__A4 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2885_ _2181_ _2163_ _2157_ mod.registers.r5\[15\] _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4512__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4624_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5234__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4555_ _1547_ _1339_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3128__I _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3506_ _2190_ _0516_ _2340_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _1317_ _1371_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2967__I _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _0368_ _0442_ _0447_ _2342_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3368_ _0374_ _0376_ _0377_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3999__S _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _1956_ _1948_ _1957_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3299_ _2404_ _0304_ _0309_ _2341_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_111_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _1345_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I io_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3446__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3461__A4 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__A1 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4174__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3921__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2877__I _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_202 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_213 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_224 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_235 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_246 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_257 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_268 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_279 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3437__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4788__I1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2670_ _2032_ _2033_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout129_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _1247_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4271_ _1252_ _1253_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3222_ _2517_ _2153_ _2519_ mod.registers.r6\[3\] _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3153_ _2414_ _2416_ _2417_ _2419_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_39_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3084_ _2140_ _2145_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3428__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3411__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4928__A1 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3986_ _0961_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2937_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3286__C _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2868_ mod.instr_2\[11\] _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _1594_ mod.registers.r1\[6\] _1582_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4156__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2799_ _2106_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3903__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4538_ _1204_ _2339_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4469_ mod.pc0\[13\] _1319_ _1471_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_104_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3419__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4417__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3198__A3 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3370__A3 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3658__A1 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _0848_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4386__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _0585_ _0704_ _0564_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2722_ mod.des.des_dout\[13\] net9 _2059_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2936__A3 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__I _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2653_ _2022_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2584_ _1985_ _1422_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5372_ _0259_ net143 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4323_ _1326_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3406__I mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout118 net125 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout129 net130 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4254_ _0820_ _2464_ _0295_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3649__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4946__B _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3850__B _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3205_ mod.registers.r1\[3\] _2234_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4185_ _0741_ _1194_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout61_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ _2432_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2872__A2 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3067_ _2218_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3141__I _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4074__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3969_ _0577_ _0858_ _0859_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3337__B1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3104__A3 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ mod.pc_1\[4\] _1819_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2606__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4872_ _1581_ mod.registers.r6\[5\] _1770_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3823_ _0554_ _0830_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4359__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3754_ _0743_ _0763_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3031__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2705_ _2051_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3685_ _0693_ _0695_ _0270_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2636_ _1989_ _2012_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3334__A3 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5355_ _0242_ net73 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2567_ mod.des.des_dout\[14\] _1973_ _1974_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _2123_ _1295_ _1297_ _1316_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5286_ _0173_ net113 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4237_ _1210_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4295__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _0767_ _1176_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_95_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ _2410_ _2227_ _2233_ mod.registers.r6\[1\] _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_55_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4047__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4099_ _0803_ _1057_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4047__B2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5318__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3022__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4430__I _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3325__A3 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__S _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4286__A1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4038__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3013__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__A1 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__B2 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4340__I _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout111_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3470_ _2231_ _0389_ _0390_ mod.registers.r6\[8\] _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5140_ _0030_ net44 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5071_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ _0578_ _1031_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4515__I _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _1805_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3806_ _0719_ _0716_ _0718_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ _1571_ _1722_ _1727_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4201__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3737_ _0745_ _0746_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4250__I _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2763__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3668_ _2267_ _0678_ _2403_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3307__A3 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4504__A2 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2619_ mod.pc_1\[8\] _2002_ _2000_ _1327_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3599_ _0325_ _0562_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5338_ _0225_ net140 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5269_ _0156_ net111 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2818__A2 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__B _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5290__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4259__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2970_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3234__A2 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4640_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4734__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _1555_ _1560_ _1562_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3522_ _2268_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3453_ _0462_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4498__B2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3384_ _0393_ mod.registers.r3\[9\] _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5123_ _0013_ net40 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5115__B _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _1800_ _1912_ _1915_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5163__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ _0857_ _0946_ _1015_ _0599_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3473__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4670__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4422__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4907_ _1508_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4973__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _1609_ _1757_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4725__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ net12 _1714_ _1514_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2736__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__A1 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__B _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3216__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4413__A1 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4964__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2975__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2559__B _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3152__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5186__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3152__B2 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2750__I1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4255__I1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2953_ mod.funct3\[2\] _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2884_ _2181_ _2172_ _2177_ mod.registers.r6\[15\] _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4623_ _1604_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4554_ _1527_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3505_ _0513_ _0514_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4485_ _2123_ _1324_ _1486_ _1487_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_fanout91_I net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ _0443_ _0444_ _0445_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ _2180_ _0375_ _2156_ mod.registers.r5\[9\] _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4891__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ mod.des.des_dout\[7\] _1951_ _1952_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3298_ _0305_ _0306_ _0307_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_57_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5037_ mod.pc\[10\] _1844_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3446__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 net22 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_203 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_214 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_225 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_236 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2893__I mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_247 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_258 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_269 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3437__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__B1 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4814__S _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3229__I _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3373__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _1256_ _1279_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3125__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3221_ _2439_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3152_ mod.registers.r4\[1\] _2228_ _2209_ mod.registers.r2\[1\] _2224_ mod.registers.r3\[1\]
+ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3083_ mod.registers.r3\[0\] _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4625__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3428__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__B _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4928__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3985_ _0992_ _0995_ _0880_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2936_ _2231_ _2227_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3600__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3139__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5351__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ _2150_ _2163_ _2164_ mod.registers.r1\[15\] _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4606_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2798_ net8 mod.des.des_dout\[28\] _2104_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4537_ mod.valid_out3 mod.ins_ldr_3 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4468_ _1291_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3116__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3419_ _2270_ _0428_ _0429_ mod.registers.r2\[11\] _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4399_ _1398_ _1404_ _1406_ _1210_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4864__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3419__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5022__C _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__B1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3758__B _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3052__B1 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3198__A4 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4304__B1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3658__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5224__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout141_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ _0529_ _0562_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3594__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2721_ _2060_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2652_ _0820_ _1797_ _1930_ mod.instr\[8\] _1809_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5371_ _0258_ net145 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2583_ _1985_ _1395_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3897__A2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _1327_ _1328_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_87_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout108 net116 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4253_ mod.pc_2\[2\] _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout119 net120 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3649__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3204_ mod.registers.r7\[3\] _2219_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3113__A4 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4184_ _2253_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3135_ _2330_ _2289_ _2292_ mod.registers.r1\[1\] _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout54_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3066_ _2358_ _2360_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2609__B1 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4074__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3578__B _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4253__I mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3968_ _0785_ _0830_ _0833_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3585__A1 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2919_ mod.registers.r5\[15\] _2201_ _2210_ mod.registers.r2\[15\] _2216_ mod.registers.r6\[15\]
+ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_3899_ _0898_ _0909_ _0818_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2702__S _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3337__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3337__B2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__I _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4837__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5247__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2699__I0 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3576__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3500__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4338__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _1824_ _1825_ _1821_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _1570_ _1777_ _1780_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3822_ _0831_ _0832_ _0325_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4006__C _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ _0698_ _0498_ _0762_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_118_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__I _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2704_ mod.des.des_dout\[5\] net18 _2049_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3684_ _0691_ _0298_ _0326_ _0351_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3319__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ _1204_ _1808_ _2011_ mod.instr\[1\] _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3417__I _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5354_ _0241_ net76 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2566_ mod.instr\[14\] _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3334__A4 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4305_ _1298_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _0172_ net126 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4819__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4236_ _1225_ _1243_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4295__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _0358_ _1177_ _0690_ _0270_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_55_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3118_ _2410_ _2415_ _2214_ mod.registers.r5\[1\] _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4098_ _1102_ _1108_ _0777_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4047__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2991__I _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3049_ _2189_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5079__I _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3022__A3 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__B1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3325__A4 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4286__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4107__B _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3549__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout90 net93 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4210__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout104_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ mod.valid1 _1903_ _1811_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4021_ _0554_ _0617_ _0620_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3788__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ mod.ins_ldr_3 _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _1661_ _1715_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3856__B _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3805_ _0538_ _0814_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4785_ mod.registers.r4\[4\] _1723_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3736_ _0682_ _2498_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3960__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3667_ _2379_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3147__I _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2618_ _1812_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3598_ _0607_ _0608_ _0350_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4504__A3 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5337_ _0224_ net138 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5268_ _0155_ net91 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4219_ mod.instr_2\[4\] _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5199_ _0089_ net74 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3243__A3 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3951__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3057__I _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2896__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4259__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3234__A3 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ mod.registers.r1\[2\] _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3942__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _2501_ _0531_ _2277_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2800__S _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ _0461_ _0448_ _0450_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4498__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3383_ _2222_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _0012_ net52 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _1913_ _1914_ _1866_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ _0878_ _0948_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3473__A3 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _1351_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3630__B1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4837_ _2530_ _1754_ _1759_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _1512_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3933__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3719_ _0728_ _0729_ _0537_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4699_ mod.registers.r2\[4\] _1671_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__A1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3924__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4120__B _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3152__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4101__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2663__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2663__B2 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2952_ _2186_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2883_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4168__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4622_ _1262_ _1605_ _1607_ _1585_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3915__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4553_ _1534_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3391__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3504_ mod.registers.r7\[14\] _2220_ _2235_ mod.registers.r1\[14\] _0515_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4484_ _1298_ _1339_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3435_ _0397_ _0389_ _0429_ mod.registers.r6\[10\] _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5130__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3366_ _2391_ _2171_ _2176_ mod.registers.r6\[9\] _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout84_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ mod.instr\[7\] _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3297_ _2410_ _2415_ _2233_ mod.registers.r4\[5\] _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5280__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _1854_ _1901_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5087__I mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4159__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4159__B2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput23 net23 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4331__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_204 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_215 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_226 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_237 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_248 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_259 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3437__A3 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5153__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3373__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3125__A2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4322__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3220_ _2517_ _2290_ _2293_ mod.registers.r5\[3\] _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3151_ _2259_ _2425_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2884__A1 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3082_ _2266_ _2379_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2636__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3984_ _0993_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4025__B _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2866_ _2157_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4605_ _1584_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2797_ _2105_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4561__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ _1529_ _1305_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4467_ mod.pc\[13\] _1292_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3116__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3418_ _2531_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4398_ _1370_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3349_ mod.pc_2\[7\] _2301_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3419__A3 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ mod.pc\[7\] _1287_ _1321_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2627__A1 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2943__B _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3052__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3052__B2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4624__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__A2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3043__A1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ mod.des.des_dout\[12\] net8 _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2651_ _2017_ _2021_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4543__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2582_ _1853_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5370_ _0257_ net143 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3897__A3 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4321_ _1329_ _1281_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ mod.pc_2\[3\] _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3203_ mod.funct7\[0\] _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4846__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4183_ _0738_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3703__I _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3134_ _2133_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3065_ _2361_ _2362_ _2199_ mod.registers.r4\[0\] _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2609__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2609__B2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4074__A3 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3859__B _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout47_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5199__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3967_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3585__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4782__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2918_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3898_ _0899_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2989__I _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2849_ _2142_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3337__A2 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3337__B3 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _1511_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2699__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2899__I mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4354__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4870_ mod.registers.r6\[4\] _1778_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3821_ _0615_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3752_ _0498_ _0762_ _0698_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2703_ _2050_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3683_ _0325_ _0310_ _0314_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3319__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2634_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _0240_ net47 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2565_ _1972_ _1970_ _1975_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4304_ _1290_ _1308_ _1309_ _1310_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_102_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _0171_ net120 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4819__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4235_ _1244_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4166_ _0890_ _0895_ _0899_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3117_ _2212_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4097_ _0977_ _1076_ _1103_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3048_ _2343_ _2344_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3255__A1 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3007__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1869_ _1418_ _1209_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2713__S _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4507__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5214__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5364__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3343__I _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3494__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4902__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3549__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net86 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net92 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__B _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2780__I0 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _0565_ _0609_ _0623_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3485__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__A3 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3202__B _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _1657_ _1747_ _1767_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3804_ _0537_ _2308_ _2354_ _0512_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__4737__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4784_ _1566_ _1722_ _1726_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3004__A4 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3735_ _0552_ _2458_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4033__B _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3666_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3872__B _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ _2001_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3597_ _2455_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4504__A4 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5336_ _0223_ net138 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2771__I0 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _0154_ net93 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ mod.ldr_hzd\[6\] _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _0088_ net63 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2708__S _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4149_ _0761_ _0505_ _0760_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3228__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__B _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3400__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4200__I0 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__I1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2690__A2 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3234__A4 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__I _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3520_ _2275_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3451_ _0448_ _0450_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3382_ _2473_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5121_ _0011_ net51 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5052_ _1913_ _1914_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _0900_ _0802_ _0655_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2681__A2 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4743__S _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4958__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _1796_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3630__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3630__B2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__I _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4836_ _1601_ _1757_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _1521_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3718_ _2311_ _0717_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4698_ _1566_ _1670_ _1672_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2997__I _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _0541_ _2242_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3697__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__C _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _0206_ net83 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3449__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3621__I _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4177__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3860__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2951_ _2242_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2882_ _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4621_ _1586_ _1324_ _1587_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4552_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3503_ mod.registers.r4\[14\] _2229_ _2225_ mod.registers.r3\[14\] _0514_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ _0442_ _0447_ _1385_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3391__A3 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3434_ _0440_ _0389_ _0390_ mod.registers.r2\[10\] _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2726__I0 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3365_ _2149_ _0375_ _2156_ mod.registers.r1\[9\] _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _1954_ _1948_ _1955_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3296_ _2408_ _2415_ _2418_ mod.registers.r1\[5\] _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ mod.pc\[9\] _1844_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4272__I _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ mod.registers.r5\[1\] _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3906__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3616__I _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_205 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_216 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_227 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_238 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_249 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4398__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3070__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4131__B _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2708__I0 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4322__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3150_ _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2884__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3081_ _2356_ _2364_ _2371_ _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__4086__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3261__I mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3046__C1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4389__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3983_ _0913_ _0867_ _0869_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4306__B _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2934_ _2197_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2865_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4604_ _1585_ _1589_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4010__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2796_ net7 mod.des.des_dout\[27\] _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4561__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4466_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4313__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ _2470_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4397_ _1322_ _1174_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3348_ _2550_ _0267_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ _2211_ mod.registers.r3\[6\] _2359_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3419__A4 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _1863_ _1877_ _1881_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2627__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__I0 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5098__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3052__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4001__A1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5047__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4304__A2 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4068__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5120__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3043__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4791__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4640__I _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__C _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2650_ _0645_ _2015_ _2019_ mod.instr\[7\] _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_fanout127_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5270__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2581_ _1854_ _1368_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4320_ _1252_ _1253_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4251_ _0487_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3202_ _2460_ _2463_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3503__B1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4182_ _0742_ _0813_ _1137_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3133_ _2427_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4059__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3064_ _2212_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__S _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__A3 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3966_ _0629_ _0877_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2917_ _2211_ _2213_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4782__A2 _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _0900_ _0351_ _0907_ _0694_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4550__I _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2848_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3337__A3 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2779_ _2095_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4518_ _1510_ mod.rd_3\[2\] _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A1 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4222__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3785__B _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4289__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ _0614_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3751_ _0505_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4764__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2775__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2702_ mod.des.des_dout\[4\] net17 _2049_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3682_ _0691_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3319__A3 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2633_ _1929_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _0239_ net50 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2564_ mod.des.des_dout\[13\] _1973_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4303_ mod.pc\[0\] _1289_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5283_ _0170_ net117 mod.pc0\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ mod.ldr_hzd\[0\] mod.ldr_hzd\[1\] mod.ldr_hzd\[2\] mod.ldr_hzd\[3\] _1245_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_101_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4165_ _0899_ _0896_ _0751_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_28_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4973__C _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3116_ mod.registers.r7\[1\] _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _1104_ _1106_ _0881_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3589__C _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3047_ mod.registers.r7\[12\] _2220_ _2235_ mod.registers.r1\[12\] _2345_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3255__A2 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__B2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4204__B2 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ mod.pc\[4\] _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3949_ _0570_ _0953_ _0958_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2766__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4507__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3191__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3494__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3246__A2 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4746__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout70 net74 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout81 net86 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2780__I1 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3485__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4365__I _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3237__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4985__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ mod.registers.r5\[15\] _1755_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3803_ _0642_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4737__A2 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ mod.registers.r4\[3\] _1723_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ _0744_ _0676_ _0616_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3665_ _2259_ _2425_ _2447_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2616_ mod.pc_1\[7\] _1996_ _2000_ _1252_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3596_ mod.pc_2\[4\] _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3173__A1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5335_ _0222_ net137 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _0153_ net92 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4217_ _1226_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5197_ _0087_ net88 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4673__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _0706_ _0463_ _1157_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_83_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4079_ _0577_ _1009_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3228__A2 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A3 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2724__S _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2739__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3400__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5331__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2679__B _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4200__I1 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3164__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2911__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2675__B1 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2978__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4913__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4134__B _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3529__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3942__A3 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3450_ _0452_ _0455_ _0459_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3155__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3381_ _0387_ _0301_ _2407_ _0388_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_112_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2902__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5120_ _0010_ net50 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4104__B1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5051_ _1445_ _1912_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4002_ _0924_ _1012_ _0646_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2608__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4028__C _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5204__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5080__A1 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4904_ _1795_ _1798_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _0285_ _1754_ _1758_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5354__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _1658_ _1706_ _1712_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3717_ _0725_ _0726_ _0727_ _0714_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ mod.registers.r2\[3\] _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3648_ _0658_ _0654_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3579_ _2502_ _2503_ _2504_ _2505_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4894__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ _0205_ net106 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5249_ _0136_ net126 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3902__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3449__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4646__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4733__I _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3385__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4885__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4908__I _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__S _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2648__B1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3860__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__I0 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4643__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _2244_ _2246_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_90_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2881_ _2166_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4620_ _1327_ _1528_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4168__A3 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1527_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3502_ mod.registers.r5\[14\] _2201_ _2210_ mod.registers.r2\[14\] _2216_ mod.registers.r6\[14\]
+ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4482_ _2123_ _1284_ _1484_ _1485_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3391__A4 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3433_ _0393_ mod.registers.r3\[10\] _0394_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2726__I1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _2546_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ mod.des.des_dout\[6\] _1951_ _1952_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _2408_ mod.registers.r3\[5\] _2223_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4628__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _1893_ _1897_ _1899_ _1309_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2639__B1 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3300__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3169__I _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _1745_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3367__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3906__A3 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4749_ _1610_ mod.registers.r3\[8\] _1699_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3119__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2590__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3833__S _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2717__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__I _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3632__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_206 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_217 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_228 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_239 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4095__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3070__A3 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3358__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3807__I _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2581__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2708__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3542__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3080_ _2372_ _2374_ _2376_ _2377_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4086__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4881__I1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5035__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3982_ _0842_ _0866_ _0883_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3046__B1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3046__C2 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4633__I1 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2933_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2864_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3349__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4603_ _1268_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2795_ _2088_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4534_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4749__S _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4465_ _1326_ _1462_ _1469_ _1288_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3416_ _0424_ _0425_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4396_ _1399_ _1400_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_98_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3347_ _0284_ _0294_ _0297_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3278_ _2367_ _2213_ _2536_ mod.registers.r4\[6\] _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4077__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5017_ _1868_ _1882_ _1885_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__I1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3588__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4001__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3512__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4458__I mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4193__I _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__C1 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3965__C _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3537__I _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3200__B1 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2580_ _1854_ _1354_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _0405_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3201_ _2482_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3503__B2 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4181_ _1143_ _1156_ _1174_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_67_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3132_ _2428_ mod.registers.r3\[1\] _2429_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4059__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3063_ _2230_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5023__A4 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3965_ _0814_ _0972_ _0975_ _0772_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2916_ _2207_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3896_ _0901_ _0902_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3990__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2847_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2778_ net16 mod.des.des_dout\[19\] _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3742__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4517_ mod.valid_out3 mod.ins_ldr_3 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4448_ _1301_ _1451_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4278__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4379_ mod.pc\[3\] _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3733__A1 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3092__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3820__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3750_ _0465_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2701_ _2043_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3681_ _0298_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _2009_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3319__A4 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _0238_ net36 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2563_ _1508_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4302_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5282_ _0169_ net120 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3216__B _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ mod.ldr_hzd\[4\] mod.ldr_hzd\[5\] mod.ldr_hzd\[6\] mod.ldr_hzd\[7\] _1244_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4164_ _0604_ _0692_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3115_ _2218_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4095_ _0783_ _0837_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout52_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3046_ mod.registers.r5\[12\] _2201_ _2210_ mod.registers.r2\[12\] _2216_ mod.registers.r6\[12\]
+ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3255__A3 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4452__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4204__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4997_ _1866_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3948_ _0593_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3177__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5309__D _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3879_ _0367_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4510__B _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3191__A2 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4140__B2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3494__A3 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3640__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout71 net74 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3954__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3087__I mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4131__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4434__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ net12 _1312_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2996__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _0527_ _1746_ _1766_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3802_ _0765_ _0773_ _0775_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4782_ _1560_ _1722_ _1725_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3733_ _2452_ _2454_ _2458_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3664_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2615_ _1931_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3595_ _0604_ _0563_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3173__A2 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4370__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5334_ _0221_ net135 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ _0152_ net92 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4122__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4216_ mod.instr_2\[3\] _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5196_ _0086_ net71 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4147_ _0937_ _0504_ _0933_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ _1008_ _0956_ _0582_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3029_ _2324_ _2326_ _2295_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4291__I _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3936__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3400__A3 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4200__I2 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3164__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2911__A2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4113__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__I _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2675__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2675__B2 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3927__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4150__B _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout102_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4352__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _2231_ _0389_ _0390_ mod.registers.r6\[9\] _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2902__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4104__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1890_ _1898_ _1905_ _1909_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4001_ _0575_ _0921_ _0885_ _1007_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__I _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2666__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2666__B2 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4407__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4903_ mod.valid0 _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3091__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2624__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4834_ _1593_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3918__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ mod.registers.r3\[15\] _1707_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4979__C _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3716_ _2313_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4591__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _1665_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3647_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4343__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3578_ _0581_ _0588_ _0550_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4995__B _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ _0204_ net103 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5248_ _0135_ net127 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3190__I _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5179_ _0069_ net68 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5179__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3082__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3909__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4582__A1 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3385__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5066__B _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4334__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4885__A2 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4637__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__I mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2648__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2648__B2 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4924__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5062__A2 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__I1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _2150_ _2172_ _2177_ mod.registers.r2\[15\] _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4573__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3501_ _0492_ _0508_ _0511_ _2313_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_7_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4481_ _0392_ _0403_ _1296_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4325__A1 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3432_ _0397_ _0400_ _0429_ mod.registers.r4\[10\] _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3363_ mod.registers.r7\[9\] _2515_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5102_ mod.instr\[6\] _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3294_ mod.registers.r7\[5\] _2413_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5033_ _1891_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2639__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2639__B2 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__B _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3367__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _1702_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3185__I _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__D _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3119__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_207 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_218 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_229 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4095__A3 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2973__B mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3070__A4 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3358__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2884__A4 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3294__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3046__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3981_ _0636_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3046__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2932_ mod.instr_2\[14\] _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2863_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3349__A2 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _1213_ _2247_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4546__B2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2794_ _2103_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4010__A3 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4533_ _1299_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4464_ _1326_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4849__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4829__I _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3415_ mod.registers.r7\[11\] _2219_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4395_ _1401_ _1377_ _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3521__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout82_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _0271_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3277_ _0285_ _2467_ _0286_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ mod.pc\[6\] _1883_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3285__A1 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4564__I _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3588__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3908__I _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5367__CLK net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3512__A2 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3276__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3818__I _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3200__A1 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3200__B2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3200_ mod.pc_2\[2\] _2483_ _2490_ _2497_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__3503__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4700__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _1179_ _1182_ _1183_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_3131_ _2144_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3062_ _2221_ mod.registers.r3\[0\] _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ _0973_ _0974_ _0643_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2915_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3895_ _0747_ _0903_ _0904_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2632__I _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2846_ mod.instr_2\[10\] _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3990__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2777_ _2089_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3742__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4516_ mod.instr_2\[5\] _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4447_ _1300_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _1356_ _1368_ _1383_ _1384_ _1386_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ mod.registers.r2\[4\] _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3258__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2743__S _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3430__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3733__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3249__A1 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3264__A4 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3421__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout132_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _2048_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3680_ _0284_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2631_ _2128_ _1797_ _1930_ mod.instr\[0\] _1809_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _0237_ net65 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2562_ _1923_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _1244_ _1245_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4379__I mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _0168_ net122 mod.pc0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4232_ _1205_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4163_ _1161_ _1163_ _1171_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3114_ _2405_ _2407_ _2409_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4094_ _0621_ _0579_ _2403_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3045_ mod.registers.r4\[12\] _2229_ _2225_ mod.registers.r3\[12\] _2343_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5003__I mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout45_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ _1859_ _1861_ _1863_ _1865_ _1867_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3947_ _0955_ _0957_ _0804_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3458__I mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3963__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3878_ _0816_ _0819_ _0823_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ mod.instr_2\[0\] _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3191__A3 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3126__C _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4140__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3651__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout61 net66 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout72 net73 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout83 net85 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4203__I0 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3706__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4199__I _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4131__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3890__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _1651_ _1743_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2996__A3 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3801_ _0798_ _0800_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_33_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4781_ mod.registers.r4\[2\] _1723_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3732_ _0643_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _0673_ _0354_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2910__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2614_ _1999_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3594_ _0361_ _0565_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3227__B _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5333_ _0220_ net139 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3173__A3 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5264_ _0151_ net89 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4215_ _2421_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _0085_ net77 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4146_ _0505_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__B _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3881__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2684__A2 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4077_ _0549_ _0784_ _0786_ _0630_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__B _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3028_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2987__A3 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1848_ _1843_ _1852_ _1847_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3936__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3400__A4 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2747__I0 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4200__I3 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2911__A3 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2675__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3624__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3098__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__I1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2730__I _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__S _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4352__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4657__I _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _0882_ _1010_ _0957_ _0878_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_78_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2666__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3091__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _1742_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3918__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4764_ _0519_ _1690_ _1711_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4040__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3715_ _0705_ _0712_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4591__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _1663_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3646_ mod.funct3\[0\] _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5250__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3577_ _0584_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _0203_ net112 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5247_ _0134_ net126 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _0068_ net67 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _0727_ _2353_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3606__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3082__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3646__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4426__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5273__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4573__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ _0509_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4480_ _2118_ _1305_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3431_ _0438_ _0301_ _0439_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4325__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _0363_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _1950_ _1948_ _1953_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3293_ _0300_ _0301_ _2407_ _0302_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _1892_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2639__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__I mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _1742_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4013__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4747_ _1602_ mod.registers.r3\[7\] _1699_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3367__A3 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3466__I _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4678_ mod.des.des_dout\[33\] _1538_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3119__A3 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _2243_ _2128_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput27 net27 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_208 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_219 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5146__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5296__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4004__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3294__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3980_ _0509_ _0659_ _0990_ _0656_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3046__A2 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2931_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2862_ mod.instr_2\[10\] _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ _1586_ _1478_ _1587_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2793_ net6 mod.des.des_dout\[26\] _2099_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4532_ _1523_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4463_ _1437_ _1463_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3414_ _2270_ mod.registers.r3\[11\] _0394_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _1373_ _1374_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5169__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3345_ _2500_ _2529_ _0353_ _0355_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout75_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3276_ mod.registers.r7\[6\] _2365_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__I0 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5015_ _1801_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4482__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3037__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4234__A1 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4785__A2 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__I _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3276__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4225__A1 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__B2 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4776__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3200__A2 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5311__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ _2139_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4665__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3061_ _2222_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3963_ _0969_ _0703_ _0713_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2914_ _2204_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3894_ _0683_ _0619_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2845_ mod.instr_2\[9\] _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2776_ _1539_ _2090_ _2093_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4515_ _1509_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4446_ _0774_ _1020_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _0342_ _0347_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3328_ mod.registers.r5\[4\] _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4575__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3259_ _0268_ _2541_ _2544_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_100_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3258__A2 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4207__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3430__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3194__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4686__S _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3497__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4694__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4446__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2733__I _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3421__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2630_ _2008_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout125_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2561_ mod.instr\[13\] _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4300_ _1225_ _1243_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5280_ _0167_ net120 mod.pc0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _1237_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4162_ _1172_ _1159_ _1160_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3113_ _2410_ _2362_ _2199_ mod.registers.r4\[1\] _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2908__I mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4093_ _0602_ _0836_ _0827_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4437__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5207__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3044_ _2341_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout38_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5357__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4995_ mod.pc\[3\] _1866_ _1509_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3946_ _0782_ _0956_ _0783_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3877_ _0856_ _0876_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2828_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4912__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2759_ _1631_ _2081_ _2083_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3191__A4 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _1412_ _1413_ _1422_ _0001_ _1435_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__4676__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4428__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3100__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2754__S _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5069__C _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout40 net45 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout51 net53 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4600__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout62 net64 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout73 net74 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2611__B1 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4903__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4667__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3890__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3987__C _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3642__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3559__I _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2996__A4 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3800_ _0496_ _0802_ _0574_ _0803_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4780_ _1551_ _1722_ _1724_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _0547_ _0667_ _0672_ _0735_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3662_ _0591_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2613_ mod.pc_1\[6\] _1996_ _1994_ _1254_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3593_ _0283_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _0219_ net139 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3173__A4 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _0150_ net89 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4214_ _1212_ _1215_ _1223_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5194_ _0084_ net77 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3243__B _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3330__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2638__I _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4145_ _1149_ _1152_ _1154_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_28_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _2262_ _1085_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3027_ _2151_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2987__A4 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _1850_ _1851_ _1319_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3397__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3929_ _0689_ _0697_ _0700_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4346__B1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3321__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3624__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3379__I _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3388__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3927__A3 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3560__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3842__I _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3312__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__S _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4901_ _1350_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _0300_ _1754_ _1756_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _1652_ _1691_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4040__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2921__I _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _0723_ _0724_ _0701_ _0699_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4694_ _1560_ _1666_ _1669_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3645_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4879__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3576_ _0585_ _0570_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4343__A3 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _0202_ net109 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5246_ _0133_ net123 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5177_ _0067_ net67 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ _0727_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__B _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ _1003_ _0879_ _1067_ _1068_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4031__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3845__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4022__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__A1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2584__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _0440_ _0398_ _2418_ mod.registers.r1\[10\] _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3361_ _0367_ _0371_ _0357_ _0299_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3572__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2887__A3 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ mod.des.des_dout\[5\] _1951_ _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3292_ _2361_ _2227_ _2199_ mod.registers.r6\[5\] _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ mod.pc\[9\] _1346_ _1380_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3836__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2916__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _1744_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4746_ _0279_ _1690_ _1701_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4677_ _1538_ _1654_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3119__A4 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628_ mod.funct3\[2\] _2245_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3559_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_209 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5229_ _0116_ net100 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A1 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4252__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2561__I mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3606__B _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3341__B _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__I mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__C _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2930_ _2221_ _2227_ _2214_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3567__I _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4172__B _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ mod.registers.r3\[15\] _2147_ _2158_ mod.registers.r4\[15\] _2159_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_30_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4600_ _1254_ _1528_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2792_ _2102_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3754__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4531_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4462_ _1465_ _1441_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3413_ _0423_ _2348_ _0422_ mod.registers.r4\[11\] _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4393_ mod.pc_2\[9\] _1374_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3344_ _2507_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ _2269_ _2474_ _2475_ mod.registers.r1\[6\] _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__I1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _1864_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout68_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__C _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3037__A3 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__I _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3745__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _1688_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4170__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4257__B _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A2 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__A4 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3984__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3387__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ _2193_ _2196_ _2357_ mod.registers.r2\[0\] _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4167__B _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ _0725_ _0726_ _0511_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3975__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2913_ _2192_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3893_ _0673_ _0622_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2844_ _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5136__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2775_ net15 _2090_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4514_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2950__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4445_ _1277_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5286__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4152__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4376_ _2117_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__I _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3327_ mod.pc_2\[4\] _2135_ _0333_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ _2541_ _2544_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4792__S _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3189_ mod.registers.r7\[2\] _2437_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4207__A2 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3430__A3 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3194__A2 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4518__I0 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4694__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A2 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3421__A3 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4382__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ _1969_ _1970_ _1971_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ _1238_ _1239_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _0821_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3112_ _2230_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4092_ _0669_ _1034_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4437__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3043_ _2257_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2999__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _1864_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3945_ _0386_ _0497_ _2380_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3876_ _0880_ _0886_ _0646_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2827_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3755__I _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4373__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2758_ mod.registers.r7\[11\] _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2689_ _2040_ _2039_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4125__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4428_ _1423_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4359_ mod.pc0\[2\] _1249_ _1363_ _1290_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_101_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4428__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5301__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout41 net43 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout63 net64 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2611__B2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout96 net97 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4203__I2 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4116__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__A2 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4419__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _0739_ _0740_ _0645_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3661_ _0545_ _0546_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2612_ _1998_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3592_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _0218_ net135 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ _0149_ net92 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3524__B _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4213_ _1205_ _0639_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2669__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5193_ _0083_ net80 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2669__B2 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3330__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4144_ _0727_ _0824_ _1141_ _0822_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4075_ _1062_ _2500_ _1063_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout50_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3026_ _2286_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2654__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _1845_ _1849_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3928_ _0760_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ _0779_ _0826_ _0495_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4346__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3944__I1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2829__I mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3321__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4585__A1 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4888__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4159__C _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _1795_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _1580_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4576__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1646_ _1706_ _1710_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _0690_ _0696_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4693_ mod.registers.r2\[2\] _1667_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3644_ _0652_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4879__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3575_ _2307_ _0570_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5314_ _0201_ net85 mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout98_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _0132_ net127 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3303__A2 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _0066_ net58 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _0509_ _0973_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _0901_ _0902_ _0906_ _0669_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_44_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4803__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ _2306_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2814__A1 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4567__A1 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3614__I0 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4319__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4774__I _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5047__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3230__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _0326_ _0327_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ mod.registers.r2\[5\] _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5030_ _1895_ _1896_ _1841_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3297__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2932__I mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _1660_ mod.registers.r5\[0\] _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4745_ _1593_ _1691_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ _1400_ _1590_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3627_ _0584_ _0580_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3763__I _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput29 net29 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4721__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3558_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3489_ _0495_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5228_ _0115_ net100 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5159_ _0049_ net48 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3003__I _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5192__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4712__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3279__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3451__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4453__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2860_ _2150_ _2154_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_fanout148_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2791_ net5 mod.des.des_dout\[25\] _2099_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4679__I _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4461_ _1437_ _1464_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3583__I mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3506__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3412_ _2203_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4392_ _2244_ _0531_ _2277_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _2525_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3274_ mod.registers.r5\[6\] _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3532__B _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2927__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5013_ _1878_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3037__A4 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4234__A3 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3993__A2 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4728_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4942__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4659_ _1552_ _1639_ _1640_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2837__I _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2572__I mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3736__A2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5110__A1 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4167__C _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3961_ _0970_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3424__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2912_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3975__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3892_ _0564_ _2403_ _0744_ _2459_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2843_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4911__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2774_ _2092_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4513_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4202__I _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3246__C _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4444_ _1258_ _1259_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2950__A3 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4375_ _2122_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout80_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ _2390_ _0334_ _0335_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3262__B _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2657__I _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3257_ mod.pc_2\[7\] _2390_ _2550_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3188_ _2428_ mod.registers.r3\[2\] _2429_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3488__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3415__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3430__A4 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4915__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3437__B _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3194__A3 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4143__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3249__A4 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3957__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3421__A4 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4206__I0 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4382__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4160_ _0761_ _0824_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3111_ _2408_ mod.registers.r3\[1\] _2223_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _0630_ _1046_ _1049_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3042_ mod.funct7\[2\] _2239_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2999__A3 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3944_ _0954_ _0781_ _0553_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4070__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3875_ _0882_ _0884_ _0885_ _0766_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2940__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2826_ mod.instr_2\[2\] _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5253__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4373__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2757_ _2064_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2688_ _1230_ _1227_ _2039_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4125__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4867__I _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4427_ _1425_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4358_ _1364_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4088__B _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2687__A2 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3309_ _2383_ _2325_ _2175_ mod.registers.r6\[5\] _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _1213_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3636__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3720__B _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3100__A3 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3011__I _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout42 net43 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout53 net60 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout75 net76 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout86 net87 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net134 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4116__A2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__I _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3875__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3875__B2 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3627__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5126__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5276__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout130_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3660_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2611_ mod.pc_1\[5\] _1996_ _1994_ _1257_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3591_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _0217_ net139 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4107__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5261_ _0148_ net93 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3166__I0 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4212_ _0423_ _1217_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3524__C _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5192_ _0082_ net54 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2669__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ _2312_ _0654_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3330__A3 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4074_ _2528_ _0749_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2935__I _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ mod.registers.r6\[12\] _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_190 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout43_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4043__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4976_ _1845_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3766__I _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ _0933_ _0937_ _0504_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3858_ _0621_ _0829_ _2338_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4346__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2809_ mod.des.des_dout\[33\] net14 _2110_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3789_ _0705_ _0656_ _0659_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__I _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3857__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5149__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3321__A3 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3609__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3450__B _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2845__I mod.instr_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4282__A1 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5299__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4034__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4585__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3545__B1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__B _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4273__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4830_ _1742_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4761_ mod.registers.r3\[13\] _1707_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3712_ _0675_ _0685_ _0688_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _1551_ _1666_ _1668_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3643_ _2252_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _2337_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5313_ _0200_ net82 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5244_ _0131_ net128 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _0065_ net48 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4500__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _0889_ _0932_ _0965_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_28_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2665__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _0675_ _0685_ _0687_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4264__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4085__C _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3008_ mod.pc_2\[13\] _2136_ _2298_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__B2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4959_ mod.pc\[11\] _1823_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2578__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4319__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__A3 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2575__I mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4007__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4730__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2741__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3290_ _2466_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_124_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3297__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__C _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3049__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3206__C1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4205__I _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _1700_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4675_ _1556_ _1504_ _1605_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2980__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3626_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3557_ _2380_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4721__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3488_ _0436_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5227_ _0114_ net123 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3288__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ _0048_ net37 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109_ _0540_ _0919_ _0791_ _0602_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4237__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _1943_ _1937_ _1944_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5337__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4712__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3771__I0 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3903__B _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3279__A2 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4228__A1 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__B2 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A2 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2790_ _2101_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4400__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2962__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _1436_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3411_ _2531_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4703__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ mod.pc_2\[10\] _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3911__B1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3342_ _0271_ _0299_ _0328_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4909__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4695__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3273_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A1 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5012_ _1880_ _1210_ _1480_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__I0 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__B1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__A3 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2988_ mod.instr_2\[11\] _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4727_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4658_ mod.registers.r1\[12\] _1526_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _0619_ _0568_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4589_ _1547_ _1452_ _1576_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2853__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A1 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2944__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4697__A1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3633__B _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ _0492_ _0508_ _0714_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2911_ _2203_ _2205_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3891_ _0892_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__A3 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2842_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3808__B _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2773_ net14 mod.des.des_dout\[17\] _2090_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ net12 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ mod.pc0\[12\] _1249_ _1446_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4374_ mod.pc0\[9\] _1369_ _1380_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_98_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3325_ _2287_ _2162_ _2392_ mod.registers.r5\[4\] _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_113_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3256_ _2432_ _0264_ _0265_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout73_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5101__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5182__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3187_ _2428_ _2484_ _2292_ mod.registers.r1\[2\] _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3663__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__B _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3415__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2623__B1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3179__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2926__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3194__A4 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3009__I _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2848__I _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3351__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3103__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2784__S _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3679__I _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4603__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2917__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4382__A3 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ _2192_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _1087_ _1094_ _1096_ _1100_ _0663_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_67_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5095__A1 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3041_ _2132_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2999__A4 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4992_ _1347_ _1312_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3943_ _2186_ _0568_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4070__A2 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3874_ _0541_ _0878_ _0603_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2825_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2756_ _2065_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2687_ _1234_ _2041_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4426_ mod.pc0\[11\] _1318_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4125__A3 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3333__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__I _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ mod.pc\[2\] _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3308_ _0315_ _0316_ _0317_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4288_ _2126_ _2128_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3239_ _2269_ _2422_ _2536_ mod.registers.r2\[7\] _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3636__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3100__A4 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__B _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout43 net45 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net56 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout76 net96 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout87 net95 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net102 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3947__I0 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3324__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3627__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4824__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4052__A2 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__A1 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2610_ _1997_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ _2462_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3563__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ _0147_ net91 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3166__I1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4211_ _1218_ _1219_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5191_ _0081_ net56 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4142_ _0737_ _2311_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3330__A4 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5068__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _0681_ _0674_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3024_ _2314_ _2317_ _2320_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_55_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_180 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_191 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3112__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5220__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout36_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4975_ _1848_ _1342_ _1320_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3926_ _0356_ _0373_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3857_ _0555_ _0866_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5370__CLK net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2808_ _1648_ _2110_ _2111_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3788_ _0704_ _0499_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4878__I _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2739_ mod.registers.r7\[3\] _2069_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4409_ _1172_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3321__A4 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3609__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__A4 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4989__S _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3545__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3545__B2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4273__A2 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _1639_ _1706_ _1709_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4191__C _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3711_ _0536_ _0720_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4691_ mod.registers.r2\[1\] _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ _0595_ _2260_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3536__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__B _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3573_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5312_ _0199_ net83 mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5243_ _0130_ net129 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3107__I mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5174_ _0064_ net36 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2946__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4125_ _0976_ _0999_ _1020_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4056_ _2526_ _1064_ _1066_ _0902_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__4264__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ _2301_ _2302_ _2303_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__A2 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _1396_ _1836_ _1835_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3775__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2578__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3909_ _0634_ _0919_ _0641_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4889_ mod.registers.r6\[13\] _1784_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3527__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5266__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__B _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2856__I _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4007__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3297__A3 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4981__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3597__I _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _1522_ _1716_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3206__B1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__C2 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3757__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ _1581_ mod.registers.r3\[5\] _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2804__I0 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4674_ _0522_ _1525_ _1653_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3625_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4221__I _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4182__A1 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3556_ _0556_ _0563_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3487_ _0497_ _0448_ _0450_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5226_ _0113_ net118 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4377__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _0047_ net37 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _0825_ _0833_ _0913_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ mod.des.des_dout\[2\] _1940_ _1941_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input16_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4237__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4039_ _0959_ _1046_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5001__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3920__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2787__S _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3771__I1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3279__A3 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3684__B1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3210__I mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4400__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2962__A2 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3410_ _0409_ _2461_ _0414_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4390_ _1370_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3911__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2697__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__B2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3341_ _0338_ _0349_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ _0273_ _0278_ _0282_ _2134_ mod.pc_2\[6\] _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ mod.pc\[6\] _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3978__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__I1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2650__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2987_ _2142_ _2163_ _2157_ mod.registers.r1\[13\] _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4726_ _1515_ _1517_ _1522_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4155__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ _2527_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4588_ _1257_ _1544_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3539_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5209_ _0099_ net88 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5304__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3969__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3433__A3 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4394__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2944__A2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2880__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__B1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3424__A3 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4621__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2910_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3890_ _0592_ _0622_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2841_ _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3188__A2 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2772_ _2091_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4511_ _1501_ _1505_ _1506_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4137__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _1291_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ _1364_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3360__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3324_ _2141_ mod.registers.r3\[4\] _2429_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3255_ _2330_ mod.registers.r3\[7\] _2145_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3115__I _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout66_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3186_ _2161_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2954__I _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__A1 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2623__B2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3179__A2 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__A3 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2926__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4709_ _1665_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4128__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3734__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3351__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3025__I mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2864__I _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__B _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3695__I _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4206__I2 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2917__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4119__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3040_ _2337_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3942_ _0583_ _0641_ _0791_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3819__B _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3873_ _0578_ _0866_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4358__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2824_ mod.des.des_counter\[1\] _0000_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2755_ _2080_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3030__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2686_ _2042_ _2041_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2949__I _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _1398_ _1426_ _1431_ _1346_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3333__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _1247_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3307_ _2493_ mod.registers.r3\[5\] _2145_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _2118_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3238_ _2198_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3169_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2695__I1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout44 net45 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout66 net97 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4349__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout77 net79 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout88 net89 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout99 net102 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3947__I1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2859__I _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3324__A2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3088__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2835__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2599__B1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3260__A1 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3012__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3563__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4210_ mod.ldr_hzd\[7\] _0394_ _1220_ mod.ldr_hzd\[6\] _2270_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5190_ _0080_ net39 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4141_ _0778_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4072_ _0733_ _1070_ _1078_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_83_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3023_ mod.registers.r5\[12\] _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_170 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_181 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_192 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ mod.pc\[1\] _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3925_ _0934_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _0831_ _0832_ _2306_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2807_ net13 _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ _0778_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2738_ _1559_ _2068_ _2071_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2669_ _0423_ _2030_ _2027_ mod.instr\[14\] _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3306__A2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ _1260_ _1261_ _1414_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3857__A3 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4339_ mod.pc0\[1\] _1313_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3490__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5195__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3545__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2589__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4309__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3213__I mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2808__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3481__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _0544_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ _1665_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3641_ _0312_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3572_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _0198_ net90 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5242_ _0129_ net129 mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _0063_ net36 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ _1039_ _1045_ _1061_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4219__I mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4055_ _0745_ _0746_ _1065_ _1063_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3123__I mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3006_ _2142_ mod.registers.r3\[13\] _2146_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3472__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4957_ mod.pc_1\[10\] _1833_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3775__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3908_ _0793_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4888_ _1638_ _1777_ _1789_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2983__B1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3839_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3793__I _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4488__B1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3033__I _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3463__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4963__A1 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5210__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3297__A4 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5360__CLK net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _1658_ _1735_ _1741_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__I0 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__B1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__B2 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _1689_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4954__A1 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2804__I1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4673_ _1582_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3624_ _0634_ _0548_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3555_ _0565_ _0503_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4182__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3486_ _0461_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout96_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _0112_ net119 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _0046_ net41 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ _0836_ _0827_ _0842_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5087_ mod.instr\[2\] _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _0949_ _1047_ _1048_ _0877_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3445__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2692__I _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3996__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4796__I1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4412__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3028__I _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3381__B1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3684__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__B2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2731__I0 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3987__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3739__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4936__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3340_ _2266_ _0350_ _0348_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4478__B _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2777__I _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3271_ _0279_ _2382_ _0280_ _0281_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _1873_ _1843_ _1879_ _1847_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__I0 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4925__C _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3978__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4927__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2986_ mod.registers.r7\[13\] _2169_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2938__B1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2789__I0 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4725_ _1658_ _1667_ _1687_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ mod.des.des_dout\[30\] _1626_ _1635_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_107_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3607_ _0616_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4155__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _1533_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3538_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3469_ _0467_ _0301_ _2407_ _0478_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_88_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__I _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5208_ _0098_ net47 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5139_ _0029_ net44 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5012__B _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3969__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2798__S _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3981__I _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3914__C _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3657__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5129__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3121__A3 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2880__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__I mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5279__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2840_ mod.instr_2\[11\] _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout146_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__A3 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2771_ net13 mod.des.des_dout\[16\] _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4510_ _2412_ _2420_ _1298_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4137__A2 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ mod.pc\[12\] _1292_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4372_ mod.pc\[9\] _1365_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3323_ _2287_ _2394_ _2396_ mod.registers.r6\[4\] _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3254_ _2330_ _2435_ _2426_ mod.registers.r2\[7\] _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3648__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4936__B _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3185_ _2432_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout59_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4999__I1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3179__A3 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2969_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _1678_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4897__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _1619_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3351__A3 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3041__I _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4119__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3327__B1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4475__C _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4990_ _1845_ _1849_ _1856_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3941_ _0808_ _0946_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3872_ _0831_ _0832_ _0790_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2823_ _2121_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4358__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2754_ _1624_ mod.registers.r7\[10\] _2077_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3030__A2 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2685_ _1230_ _1232_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _1370_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ _1288_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3333__A3 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3306_ _2493_ _2325_ _2395_ mod.registers.r2\[5\] _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4286_ _2472_ _2480_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2965__I _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3237_ mod.registers.r7\[7\] _2365_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3168_ _2202_ _2204_ _2206_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3099_ _2391_ _2394_ _2396_ mod.registers.r6\[0\] _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout45 net46 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout56 net59 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout67 net69 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4349__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout78 net79 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout89 net94 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3324__A3 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2875__I mod.instr_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2835__A2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2599__B2 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3260__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3012__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4140_ _0637_ _0955_ _1150_ _0898_ _0880_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_110_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4071_ _2262_ _1003_ _1067_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_68_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3022_ _2318_ _2319_ _2292_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_55_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_160 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_171 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_182 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_193 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4028__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _1842_ _1843_ _1846_ _1847_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3924_ _0476_ _0486_ _0488_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3251__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3855_ _0789_ _0829_ _0529_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2806_ mod.des.des_counter\[2\] _2122_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3786_ _0788_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2737_ mod.registers.r7\[2\] _2069_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4240__I _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2762__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2668_ _1988_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3306__A3 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4407_ _1263_ _1273_ _1274_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4503__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2599_ mod.pc_1\[0\] _1990_ _1933_ mod.pc_2\[0\] _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4269_ mod.pc_2\[6\] _1255_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5071__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4616__S _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4019__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3490__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4814__I0 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3617__I1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3475__B _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4258__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _2462_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5310_ _0197_ net88 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _0128_ net128 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5172_ _0062_ net43 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ _1083_ _1101_ _1115_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__I mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4054_ _0747_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 io_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3005_ _2142_ _2172_ _2177_ mod.registers.r2\[13\] _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3472__A2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _1381_ _1834_ _1835_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3907_ _0916_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ mod.registers.r6\[12\] _1778_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2983__B2 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3838_ _0657_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4724__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ _2306_ _0779_ _0615_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2735__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4488__B2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3160__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3463__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__B1 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3917__C _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4715__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3151__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4100__B1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ mod.registers.r4\[15\] _1736_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__A2 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__B2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4254__I1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _1571_ _1693_ _1698_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__A2 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4706__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3623_ _2507_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3554_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3485_ _0495_ _0436_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _0111_ net123 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout89_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _0045_ net40 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3134__I _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4890__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ _0806_ _0912_ _0914_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5086_ _1939_ _1937_ _1942_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ _0913_ _0858_ _0861_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3445__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4939_ mod.pc_1\[3\] _1819_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3044__I _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2731__I1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2883__I _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2798__I1 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__I _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3372__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3270_ mod.registers.r2\[6\] _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3889__I _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2635__B1 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2985_ _2189_ _2282_ _2241_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2938__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2789__I1 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2938__B2 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ mod.registers.r2\[15\] _1675_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4655_ _1535_ _1636_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3606_ _2268_ _0579_ _2448_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4586_ _1533_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3363__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3537_ _2482_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5104__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3468_ mod.registers.r7\[8\] _2413_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _0097_ net47 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3399_ mod.registers.r7\[11\] _2515_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4863__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2713__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _0028_ net68 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5069_ _1500_ _1927_ _1928_ _1853_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3969__A3 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4918__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5040__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5350__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3354__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2704__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__A4 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3409__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3658__B _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout139_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2770_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3393__B _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3345__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _1321_ _1372_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_125_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ _0329_ _0330_ _0331_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3253_ _2324_ _2319_ _2426_ mod.registers.r4\[7\] _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3648__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3184_ _2258_ _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5223__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__B _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__A1 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4243__I mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2968_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4707_ _1602_ mod.registers.r2\[7\] _1663_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2899_ mod.instr_2\[12\] _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4638_ _0449_ _1576_ _1621_ _1585_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4569_ _1524_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5074__I _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4836__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3272__B1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3024__B1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3575__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3327__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3327__B2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4102__B _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4827__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3940_ _0947_ _0948_ _0950_ _0636_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3871_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5004__A1 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2822_ mod.des.des_counter\[2\] _2114_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__I mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2753_ _2079_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2684_ _2040_ _2041_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3318__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4423_ _2238_ _0409_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3407__I mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3333__A4 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3851__B _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ mod.registers.r7\[5\] _2167_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4285_ _2117_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3570__C _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout71_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3236_ _2530_ _2467_ _2532_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4294__A2 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3167_ mod.registers.r5\[2\] _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3098_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout46 net61 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout57 net59 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout68 net69 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout79 net87 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4701__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3309__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5269__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2599__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3720__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4070_ _0875_ _0987_ _1079_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3021_ _2160_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_161 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_172 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_183 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_194 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _1805_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3787__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3923_ _0503_ _0489_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3854_ _0860_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2805_ _2109_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3785_ _0766_ _0792_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ _1550_ _2068_ _2070_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2667_ _2025_ _2031_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4406_ _0288_ _0293_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2598_ _1812_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2976__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4268_ _1258_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3219_ _2324_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4199_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4814__I1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__A3 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4258__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4606__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout121_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4341__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3570_ _0530_ _0575_ _0578_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3941__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5240_ _0127_ net128 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5171_ _0061_ net38 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4122_ _1123_ _1127_ _1129_ _1132_ _0663_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ _1062_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3457__B1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 io_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3004_ _2288_ _2163_ _2177_ mod.registers.r4\[13\] _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3472__A3 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4516__I mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3209__B1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2680__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _1794_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3906_ _0783_ _0830_ _0859_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4886_ _1631_ _1777_ _1788_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3837_ _0594_ mod.funct3\[1\] _2260_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4251__I _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3768_ _0614_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ _2043_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3699_ _0707_ _0708_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4488__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ _0256_ net136 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5082__I mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3160__A2 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5307__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3463__A3 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__B _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__B2 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4161__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3923__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3933__C _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3151__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4100__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4100__B2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__B _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ mod.registers.r3\[4\] _1694_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ _1648_ _1626_ _1649_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4167__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3622_ _0631_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3553_ _0561_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3484_ _0493_ _0416_ _0419_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5223_ _0110_ net114 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3142__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ _0044_ net49 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4105_ _0626_ _0553_ _0866_ _0883_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ mod.des.des_dout\[1\] _1940_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4036_ _0863_ _0870_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__A3 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4246__I mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3150__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ mod.pc\[3\] _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4869_ _1565_ _1777_ _1779_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4158__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3905__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3381__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4149__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__B1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__B2 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2984_ _2279_ _2280_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _0526_ _1666_ _1686_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2938__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3060__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4015__B _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _1253_ _1599_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3605_ _0614_ _0615_ _2402_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4585_ mod.des.des_dout\[23\] _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3536_ _2264_ _0545_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4560__A1 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3363__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ mod.registers.r2\[8\] _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5206_ _0096_ net71 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3398_ mod.pc_2\[11\] _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5137_ _0027_ net68 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ net19 _1500_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input14_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ _0631_ _0958_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4091__A3 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3051__A1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3764__B _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4000__B1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3354__A2 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__A1 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2894__I _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2880__A4 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3042__A1 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4370_ _1326_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ _2287_ _2162_ _2495_ mod.registers.r4\[4\] _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ _2545_ _2547_ _2548_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__C1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3183_ _2240_ _2339_ _2464_ _2472_ _2480_ _2355_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ _2257_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4706_ _0281_ _1674_ _1677_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4781__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ _1586_ _1405_ _1587_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4399__C _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3519_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1411_ _2237_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4836__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3639__A3 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5090__I mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3603__I _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A3 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3759__B _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3272__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3272__B2 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A2 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2889__I _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3327__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_310 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3669__B _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout151_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _0592_ _0877_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5004__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2821_ _2120_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2752_ _1616_ mod.registers.r7\[9\] _2077_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2683_ _1224_ _1807_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3318__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _1399_ _1400_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A3 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4353_ _1283_ _1358_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3304_ _2286_ _2161_ _2395_ mod.registers.r4\[5\] _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ mod.pc0\[7\] _1249_ _1287_ _1290_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3235_ _2203_ _2205_ _2531_ mod.registers.r4\[7\] _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout64_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ mod.instr_2\[5\] _2361_ _2373_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5340__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3097_ _2173_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3254__A1 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout36 net38 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout47 net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout69 net75 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3999_ _1008_ _1009_ _0949_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4754__A1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3309__A2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4809__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3493__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A3 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3245__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3796__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4113__B _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3508__I mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2568__B _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3020_ _2166_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_162 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_173 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_184 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_195 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3236__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _1844_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _0408_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3251__A4 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3853_ _0554_ _0861_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4736__A1 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2804_ net11 mod.des.des_dout\[31\] _2089_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3784_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2735_ mod.registers.r7\[1\] _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3418__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2666_ _0428_ _2030_ _2027_ mod.instr\[13\] _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4405_ _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2597_ _1989_ _1474_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4336_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4249__I mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4267_ _1259_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3218_ mod.registers.r7\[3\] _2515_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3475__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4198_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2992__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3149_ _2431_ _2434_ _2443_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__A4 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5236__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3328__I mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3063__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3218__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4108__B _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3012__B _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4718__A1 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3238__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout114_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3941__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _0060_ net49 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2752__I0 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4121_ _0749_ _0670_ _1128_ _1130_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4052_ _0673_ _2525_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3457__B2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 io_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3003_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3209__B2 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4957__A1 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ mod.pc_1\[9\] _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5259__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ _0785_ _0858_ _0861_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ mod.registers.r6\[11\] _1778_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4532__I _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3836_ _0633_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3767_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _2058_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3698_ _0556_ _0404_ _0406_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2649_ _2017_ _2020_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5368_ _0255_ net136 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3696__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2743__I0 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4319_ mod.pc_2\[7\] _1253_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5299_ _0186_ net106 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3448__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3611__I _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3463__A4 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4100__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__A1 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _1374_ _1590_ _1542_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _0598_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3552_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3914__A2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3483_ _0409_ _2461_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _0109_ net110 mod.ri_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5153_ _0043_ net51 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4104_ _1109_ _1110_ _1114_ _1112_ _0663_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_57_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _1801_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _0549_ _0993_ _0994_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__A4 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3602__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ _1424_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4868_ mod.registers.r6\[3\] _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4158__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3819_ _0621_ _0829_ _0604_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4799_ _0453_ _1719_ _1734_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2711__S _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3905__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__I mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3669__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3841__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4641__I0 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__I _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2576__B _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4085__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4085__B2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2635__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4388__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2983_ mod.registers.r4\[13\] _2229_ _2235_ mod.registers.r1\[13\] _2281_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4722_ _1652_ _1679_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3060__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _1545_ _1443_ _1605_ _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3604_ _0560_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3899__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4584_ _1519_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3535_ _0544_ _0538_ _0539_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4560__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3466_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4966__B _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _0095_ net65 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3397_ _0386_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5136_ _0026_ net54 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _1224_ _0649_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4076__A1 _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4018_ _1025_ _1027_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2706__S _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4000__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__B2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3814__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4790__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3320_ mod.registers.r7\[4\] _2168_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3251_ _2318_ _2435_ _2439_ mod.registers.r6\[7\] _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__B1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3502__C2 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3182_ _2476_ _2477_ _2478_ _2479_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3805__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3281__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2966_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4705_ _1594_ _1675_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4781__A2 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2897_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _1399_ _1528_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4567_ mod.des.des_dout\[20\] _1543_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3518_ _0521_ _0524_ _0528_ _2136_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_103_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _1317_ _1443_ _1452_ _1356_ _1496_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2995__I _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3449_ mod.pc_2\[10\] _2390_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _0009_ net42 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3272__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3024__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_300 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2820_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout144_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3685__B _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2751_ _2078_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4763__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2682_ _1226_ _1227_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _1401_ _1377_ _1427_ _1402_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3318__A3 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4352_ _1359_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3303_ _2542_ _0311_ _0313_ _2265_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4283_ _1291_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3234_ _2469_ _2470_ _2531_ mod.registers.r6\[7\] _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3165_ _2462_ _2448_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3096_ _2325_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout57_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3254__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout37 net38 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout59 net60 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3006__A2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3998_ _0691_ _0366_ _0564_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4754__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2949_ _2188_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4506__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _1533_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__C _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5165__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3493__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3245__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4442__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4745__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__C _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3181__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_152 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_163 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_174 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_185 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_196 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4970_ _1842_ _1308_ _1320_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3236__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3921_ _0911_ _0926_ _0930_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_63_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4984__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2804__S _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3852_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2803_ _2108_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4736__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ _0634_ _0793_ _0641_ _2185_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2734_ _2064_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2665_ _1424_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ _2113_ mod.des.des_counter\[0\] _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2596_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4335_ mod.valid2 _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4266_ _1260_ _1261_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3217_ _2167_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3475__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4197_ _2130_ _1206_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3148_ _2444_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _2272_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2986__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2738__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5045__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3218__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__B2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3519__I _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5330__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3154__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ _2499_ _0680_ _0879_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2752__I1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4051_ _0548_ _0619_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3457__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4654__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3002_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4406__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2680__A3 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _1388_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4957__A2 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4813__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3904_ _0808_ _0912_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4884_ _1787_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3835_ _0627_ _0835_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3429__I _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3766_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3393__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ mod.des.des_dout\[11\] net7 _2054_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3697_ _0486_ _0488_ _0476_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2648_ _0738_ _2015_ _2019_ mod.instr\[6\] _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5367_ _0254_ net136 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2579_ _1984_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3696__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4893__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2743__I1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4318_ _2278_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5298_ _0185_ net106 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ mod.pc_2\[4\] _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5203__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5353__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3783__B _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3136__A1 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3439__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5117__RN _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__I0 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3620_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3551_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3482_ _0410_ _0411_ _0412_ _0413_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3127__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _0108_ net103 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5152_ _0042_ net52 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3142__A4 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4103_ _0662_ _1111_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _1924_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4627__A1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _0671_ _1041_ _1044_ _0733_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5376__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4936_ _1366_ _1822_ _1821_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3602__A2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _1769_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3818_ _2379_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4798_ _1623_ _1720_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3366__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2998__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3905__A3 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3749_ _0756_ _0757_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3118__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3669__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__B1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3841__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4641__I1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3069__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2701__I _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2580__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5249__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4609__A1 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3293__B1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3045__B1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2982_ mod.registers.r7\[13\] _2220_ _2225_ mod.registers.r3\[13\] _2280_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _1646_ _1667_ _1685_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3060__A3 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ _1464_ _1529_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3603_ _0559_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4583_ _1555_ _1571_ _1572_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3534_ _0538_ _0539_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2571__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3465_ _0468_ _0471_ _0475_ _2483_ mod.pc_2\[8\] _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__4848__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _0094_ net65 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout87_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3396_ _0404_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5135_ _0025_ net55 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5066_ _1925_ _1926_ _1841_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4017_ _0598_ _0992_ _0948_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3823__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3598__B _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A1 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _1807_ _1810_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2722__S _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3339__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4000__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4303__A3 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__B _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A1 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4116__C _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3578__A1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3042__A3 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2553__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3250_ _2179_ _2319_ _2441_ mod.registers.r5\[7\] _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3181_ mod.registers.r7\[2\] _2218_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3805__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3281__A3 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3569__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2965_ _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4704_ _0302_ _1674_ _1676_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4821__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3865__C _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2896_ mod.instr_2\[13\] _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ mod.des.des_dout\[28\] _1542_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4566_ _1556_ _1360_ _1546_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3741__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3517_ _0525_ _2510_ _0280_ _0526_ _2320_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _1412_ _0516_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3448_ _2300_ _0456_ _0457_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4297__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _2232_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _0008_ net42 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4049__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5049_ mod.pc\[12\] _1903_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2717__S _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5099__I _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3272__A3 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3980__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4288__A2 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_301 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2750_ _1610_ mod.registers.r7\[8\] _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout137_I net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3971__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2681_ _1234_ _2039_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ mod.pc_2\[10\] _1400_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3318__A4 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _1302_ _1133_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_125_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ _0312_ _2542_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4282_ mod.pc\[7\] _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3233_ _2197_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3164_ _2461_ _2425_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4816__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3095_ _2391_ _2162_ _2392_ mod.registers.r5\[0\] _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4451__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__B _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout38 net46 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net53 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3997_ _0361_ _0503_ _2380_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3006__A3 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2948_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3962__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3167__I mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4618_ mod.des.des_dout\[26\] _1573_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3309__A4 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3714__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _1519_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4410__B _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3181__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3469__B1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3484__A3 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4681__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_153 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_164 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_175 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_186 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_197 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4433__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3920_ _2264_ _0897_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3696__B _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3851_ _2267_ _0678_ _0461_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2802_ net10 mod.des.des_dout\[30\] _2104_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3782_ _0608_ _0348_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2733_ _2065_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2664_ _2025_ _2029_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4403_ _1356_ _1395_ _1409_ _1384_ _1410_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_2595_ _1793_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4334_ _2130_ _1206_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__S _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4265_ _1263_ _1273_ _1274_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4121__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3216_ _2513_ _2317_ _2483_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4196_ mod.valid2 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3475__A3 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3147_ _2257_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2683__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3078_ _2251_ _2375_ _2272_ _2208_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2986__A2 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4281__I _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2738__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5132__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4230__B _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3625__I _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2674__A1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4103__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ _0822_ _1041_ _1051_ _0646_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_84_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3001_ _2133_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3270__I mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4406__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _1335_ _1832_ _1829_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3903_ _0867_ _0869_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3090__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ _1624_ mod.registers.r6\[10\] _1772_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3834_ _0627_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__C _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3917__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3765_ _2252_ _2254_ _0596_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_118_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3393__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2716_ _2057_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3696_ _0404_ _0406_ _0556_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2647_ _1929_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5366_ _0253_ net136 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2578_ _0003_ _1315_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4893__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ mod.pc_2\[8\] _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5297_ _0184_ net117 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _1257_ _0449_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4276__I _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4179_ _0751_ _0824_ _1187_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2656__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5070__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2959__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3081__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__C _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3384__A2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4186__I _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4914__I _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3072__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5178__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _0559_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3481_ _0356_ _0373_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3127__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4324__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _0107_ net110 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ _0041_ net53 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4102_ _0821_ _0650_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ mod.instr\[1\] _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4627__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _1042_ _1043_ _0766_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3438__I0 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4935_ mod.pc_1\[2\] _1819_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4866_ _1772_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3817_ _0583_ _0825_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4797_ _1733_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3366__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3748_ _0758_ _0709_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3679_ _0269_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3175__I _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3118__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5349_ _0236_ net63 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4618__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__A1 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__B2 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3054__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__I _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3293__A1 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3293__B2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__A2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3045__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2981_ mod.registers.r5\[13\] _2201_ _2210_ mod.registers.r2\[13\] _2216_ mod.registers.r6\[13\]
+ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3045__B2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ mod.registers.r2\[13\] _1675_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3060__A4 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4651_ _1555_ _1632_ _1633_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3602_ _0603_ _0606_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4582_ mod.registers.r1\[4\] _1561_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3533_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3464_ _2134_ _0472_ _0473_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5203_ _0093_ net39 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4848__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3723__I _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3395_ _2266_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5134_ _0024_ net41 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ mod.valid1 _1806_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _0677_ _0852_ _1026_ _2449_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3284__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__A3 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4784__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4918_ mod.rd_3\[2\] _1808_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4849_ _1645_ _1747_ _1765_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3339__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4729__I _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3275__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4775__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4527__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5216__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5366__CLK net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3543__I _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__A2 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3180_ _2469_ _2474_ _2232_ mod.registers.r4\[2\] _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_66_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3266__A1 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3281__A4 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3569__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4766__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2964_ _2253_ _2254_ _2261_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ _1580_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2895_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _1618_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ _1264_ _1536_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3741__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3516_ mod.registers.r5\[14\] _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4496_ _1384_ _1426_ _1495_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4549__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3447_ _2141_ _0375_ _2156_ mod.registers.r1\[10\] _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_103_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3378_ _2470_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5117_ _0007_ _0003_ net145 mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _1868_ _1910_ _1911_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3257__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__B1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3980__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2791__I0 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__I mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_302 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4194__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4996__B2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4922__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3420__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3538__I _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3971__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2680_ _1510_ _1224_ _1813_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ _1250_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4920__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3301_ mod.funct3\[0\] _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2782__I0 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4281_ _1247_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3273__I _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3232_ mod.registers.r5\[7\] _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3487__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input4_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3163_ _2265_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3239__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3094_ _2291_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__B2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3254__A4 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4739__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout39 net40 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3996_ _0857_ _0955_ _0593_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2947_ _2240_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2878_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4617_ _1603_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _2387_ _1525_ _1541_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2773__I0 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _2123_ _1474_ _1482_ _1483_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3478__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__I _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3469__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__I _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_154 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_165 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_176 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_187 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_198 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ _0779_ _0826_ _0556_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2801_ _2107_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3781_ _0568_ _0582_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3268__I mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2732_ _2067_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2663_ _1216_ _2023_ _2027_ mod.instr\[12\] _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _0304_ _0309_ _1385_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2594_ _1987_ _1449_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4333_ _1338_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4264_ _1260_ _1261_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3215_ mod.registers.r1\[3\] _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4121__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4195_ _1196_ _1203_ _1204_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3146_ mod.pc_2\[1\] _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4048__B _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3077_ _2124_ _2127_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_54_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3979_ _0509_ _0650_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__I1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3641__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4179__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4351__A2 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3000_ _2284_ _2285_ _2294_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 io_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ mod.pc_1\[8\] _1827_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3902_ _0552_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3090__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4882_ _1786_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3833_ _0838_ _0841_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3764_ _0763_ _0764_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2715_ mod.des.des_dout\[10\] net6 _2054_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3393__A3 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3726__I _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _0462_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2646_ _2017_ _2018_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4342__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ _0252_ net135 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2577_ _1982_ _1925_ _1983_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4316_ _1301_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5296_ _0183_ net98 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4247_ _1257_ _0449_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4178_ _0270_ _0656_ _0599_ _0628_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_67_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ _2324_ _2289_ _2426_ mod.registers.r4\[1\] _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3605__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3384__A3 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4333__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3844__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3072__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout112_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ _0408_ _0437_ _0465_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_6_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3127__A3 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _0040_ net41 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4101_ _0616_ _0841_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5081_ _1935_ _1937_ _1938_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4088__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4032_ _0723_ _0724_ _0936_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__I0 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3438__I1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4934_ _1352_ _1820_ _1821_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4260__A1 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4865_ _1559_ _1773_ _1776_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3816_ _0614_ _0826_ _0354_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4012__A1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1617_ mod.registers.r4\[9\] _1728_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3747_ _0386_ _0407_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3366__A3 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3678_ _0675_ _0685_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4315__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2629_ mod.pc_1\[13\] _1813_ _1932_ mod.pc_2\[13\] _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5348_ _0235_ net62 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4287__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3405__B _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4079__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _0166_ net100 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2629__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__I0 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4306__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3315__B _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3293__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5295__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2980_ _2270_ _2275_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3045__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4650_ mod.registers.r1\[11\] _1561_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 io_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3601_ _0603_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4581_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3532_ _0541_ _2242_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3463_ _2488_ _2484_ _2495_ mod.registers.r4\[8\] _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _0092_ net89 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3394_ mod.funct7\[1\] _2332_ _2274_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _0023_ net72 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3808__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _0677_ _0801_ _0655_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4481__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3284__A2 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3036__A2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A1 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3895__B _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4917_ _1509_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4784__A2 _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ mod.registers.r5\[13\] _1755_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3186__I _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ mod.registers.r4\[1\] _1723_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5168__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3275__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4472__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3096__I _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3018__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2963_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2903__I _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4702_ _1662_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2894_ _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4633_ _1617_ mod.registers.r1\[9\] _1554_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3935__S _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _2130_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3515_ mod.registers.r2\[14\] _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5310__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _1298_ _1493_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3446_ mod.registers.r7\[10\] _2515_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3377_ mod.registers.r2\[9\] _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5116_ _1961_ _1959_ _1964_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ mod.pc\[11\] _1883_ _1884_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3257__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__B2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2768__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3193__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2791__I1 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4693__A1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_303 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__A2 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2759__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3420__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5333__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3971__A3 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3184__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3554__I _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4920__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3300_ _2372_ _2374_ _2376_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_125_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2782__I1 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _1289_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3231_ _2526_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3487__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3162_ _2380_ _2403_ _2449_ _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_94_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3093_ _2383_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3239__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4987__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__A2 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ _0898_ _1002_ _1005_ _0818_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2877_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _1602_ mod.registers.r1\[7\] _1554_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _1526_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4911__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ _0480_ _0485_ _1296_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3429_ _2473_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5356__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3402__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2764__I1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3469__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4418__A1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_155 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_166 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_177 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_188 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_199 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4154__B _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout142_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2800_ net9 mod.des.des_dout\[29\] _2104_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3780_ _0789_ _0790_ _2481_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2731_ _1660_ mod.registers.r7\[0\] _2066_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2601__B1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2662_ _2025_ _2028_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2593_ _1425_ _1433_ _1815_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4332_ _1301_ _1339_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ mod.pc_2\[3\] _1262_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5229__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3214_ _2508_ _2509_ _2510_ _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4121__A3 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4194_ _0661_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3145_ _2436_ _2438_ _2440_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3076_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _0978_ _0981_ _0983_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3396__A1 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2929_ _2195_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3148__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3922__I _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4820__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4887__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3832__I _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput8 io_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3988__B _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4950_ _1293_ _1831_ _1829_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4811__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3901_ _0863_ _0870_ _0842_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4881_ _1617_ mod.registers.r6\[9\] _1772_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3832_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3763_ _2263_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _2056_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3694_ _0704_ _0499_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2645_ _1510_ _2015_ _2011_ mod.instr\[5\] _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _0251_ net139 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2576_ mod.des.des_dout\[17\] _1936_ _1509_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3550__A1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4315_ _1251_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _0182_ net98 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4246_ mod.pc_2\[5\] _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3302__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4177_ _0690_ _0853_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3853__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3128_ _2174_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5055__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _2198_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3081__A3 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3369__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2821__I _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2592__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3652__I _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3780__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2583__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout105_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3532__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _0852_ _0679_ _1105_ _0850_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ mod.des.des_dout\[0\] _1925_ _1884_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4594__S _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ _0700_ _0689_ _0697_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3835__A2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__I1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1794_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4260__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ mod.registers.r6\[2\] _1774_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3815_ _0615_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4795_ _1732_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4012__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__I _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _0504_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3366__A4 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2574__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3677_ _0357_ _0686_ _0328_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2628_ _2007_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3118__A4 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5347_ _0234_ net82 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2559_ mod.des.des_dout\[12\] _1962_ _1963_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5278_ _0165_ net121 mod.pc0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4079__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4229_ _0661_ _0639_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4874__I1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5028__A1 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3039__B1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2752__S _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4003__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2551__I mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3762__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3382__I _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__I mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3600_ _0563_ _0609_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput11 io_in[19] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_30_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ mod.des.des_dout\[22\] _1543_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3531_ _2137_ _0540_ _2249_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2556__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2800__I0 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3462_ _2494_ mod.registers.r3\[8\] _2429_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _0091_ net78 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__B _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3393_ _2356_ _0392_ _0403_ _2342_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_69_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _0022_ net57 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _0821_ _1022_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4481__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3036__A3 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A2 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4916_ _1424_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3441__B1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4072__B _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__I mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _1638_ _1747_ _1764_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4778_ _1717_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3744__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__I0 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3729_ _0737_ _2250_ _0736_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_107_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2747__S _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3151__B _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3275__A3 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__A2 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3983__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3735__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4160__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3840__I _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5262__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3266__A3 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__S _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3996__B _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3018__A3 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2962_ _2256_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4701_ _1663_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3974__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2893_ mod.instr_2\[14\] _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4632_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3514_ mod.registers.r4\[14\] _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4494_ _1411_ _2282_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3445_ _2391_ _2171_ _2176_ mod.registers.r6\[10\] _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3376_ mod.registers.r5\[9\] _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_fanout85_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ mod.des.des_dout\[9\] _1962_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1908_ _1909_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__B _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__I _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2768__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3197__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3717__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3193__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4142__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4693__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4756__I _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3660__I _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_304 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3653__B1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3420__A3 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3184__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3771__S _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3230_ _2482_ _2527_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4133__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3161_ _2452_ _2454_ _2458_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_67_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3092_ _2299_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3239__A3 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__A2 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ _0895_ _1004_ _0643_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5158__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2945_ mod.funct7\[1\] _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2876_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__I0 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4615_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4372__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4546_ _1530_ _1535_ _1537_ _1538_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _2118_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4124__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3428_ mod.registers.r7\[10\] _2413_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4675__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3359_ _2243_ _0368_ _0369_ _2246_ _0338_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ mod.pc\[8\] _1843_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3402__A3 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3390__I _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2677__A1 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_156 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4418__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_167 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_178 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_189 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2734__I _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3929__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2601__A1 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2601__B2 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _2181_ _2023_ _2027_ mod.instr\[11\] _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3565__I _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ _1338_ _1396_ _1397_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2592_ _1987_ _1409_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _1300_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4106__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4262_ _1264_ _1265_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3213_ mod.registers.r4\[3\] _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4193_ _2246_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3144_ _2318_ _2319_ _2441_ mod.registers.r5\[1\] _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A3 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3075_ mod.funct3\[2\] _2255_ _2132_ _2239_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_54_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__I _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3977_ _0959_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3396__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2928_ mod.registers.r7\[15\] _2220_ _2225_ mod.registers.r3\[15\] _2226_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2859_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3148__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _1515_ _1518_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2819__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4820__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2554__I mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2729__I _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3311__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3075__A1 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4165__B _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3900_ _0743_ _0897_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2822__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _0469_ _1773_ _1785_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3831_ _0601_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3762_ _0767_ _0771_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2713_ mod.des.des_dout\[9\] net5 _2054_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3693_ _0421_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2644_ _1988_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _0250_ net135 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2575_ mod.instr\[17\] _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3550__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4314_ _1322_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5294_ _0181_ net98 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ _1254_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5015__I _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4176_ _1185_ _1186_ _0961_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3853__A3 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3127_ _2404_ _2412_ _2420_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_27_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3058_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3369__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4869__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3154__B _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3072__A4 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A1 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5219__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3780__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3517__C1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__CLK net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3532__A2 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _0756_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3296__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5037__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3599__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ mod.pc_1\[1\] _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _1550_ _1773_ _1775_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4548__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2922__I _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ _2309_ _0678_ _0338_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4794_ _1610_ mod.registers.r4\[8\] _1728_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3745_ _0754_ _0755_ _0700_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3220__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3676_ _0352_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2627_ mod.pc_1\[12\] _1813_ _1932_ _1464_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3523__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4720__A1 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _0233_ net82 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2558_ _1924_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _0164_ net99 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4228_ mod.ldr_hzd\[0\] _1231_ _1228_ mod.ldr_hzd\[2\] mod.instr_2\[5\] _1239_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4584__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4159_ _0778_ _1165_ _1167_ _0874_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3039__B2 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3612__B _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3817__A3 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__I0 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput12 io_in[1] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3530_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3753__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4950__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2800__I1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3461_ _2494_ _2394_ _2396_ mod.registers.r2\[8\] _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3573__I _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ _0090_ net71 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3392_ _0395_ _0396_ _0399_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _0021_ net70 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ mod.valid0 _1347_ _1811_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4013_ _1022_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A3 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _1510_ _1805_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3441__A1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4846_ mod.registers.r5\[12\] _1755_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _1718_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3744__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4941__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__I1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3728_ _2250_ _0736_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3659_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _0216_ net142 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3275__A4 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2562__I _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__A2 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4932__A1 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3499__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5113__I _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3266__A4 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2961_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3568__I _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _1571_ _1670_ _1673_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3974__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2892_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _1612_ _1615_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _1524_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3513_ _0522_ _2317_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4493_ _1460_ _1083_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3444_ _0453_ _2510_ _0280_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3375_ _0384_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _1508_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2647__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ mod.pc\[11\] _1903_ _1432_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3414__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _1743_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3193__A3 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_305 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2557__I mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3653__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4772__I _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__A4 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5108__I mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _2444_ _2455_ _2456_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__3892__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__S _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3091_ _2387_ _2316_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3239__A4 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3644__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__I _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ _1000_ _1003_ _0370_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2944_ _2190_ _2237_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2875_ mod.instr_2\[9\] _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _1596_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__I1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4545_ mod.des.des_dout\[18\] _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3580__B1 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4476_ _1290_ _1475_ _1476_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ mod.registers.r5\[10\] _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3761__I _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4675__A3 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3358_ _0342_ _0347_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2686__A2 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3289_ mod.registers.r5\[5\] _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _1883_ _1893_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input10_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4592__I _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3001__I _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3402__A4 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2840__I mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5252__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4363__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4767__I _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3874__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2677__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_157 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4418__A3 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_168 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_179 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4051__A1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3846__I _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2601__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2660_ _1929_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2591_ _1987_ _1383_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4330_ _1267_ _1269_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3581__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _1267_ _1269_ _1270_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3212_ _2384_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _0645_ _1199_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_95_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _2291_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3074_ mod.instr_2\[3\] _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5275__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3976_ _0806_ _0984_ _0985_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2927_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3756__I _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2660__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2858_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4788__S _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2789_ net4 mod.des.des_dout\[24\] _2099_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4528_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ mod.pc_2\[12\] _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3084__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2831__A2 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3847__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5148__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3311__A3 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5298__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3075__A2 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3830_ _0565_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4024__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3761_ _0662_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2586__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ _2055_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3692_ _0689_ _0697_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4327__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2643_ _1989_ _2016_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _0249_ net140 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2574_ _1980_ _1925_ _1981_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4313_ _1045_ _1061_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5293_ _0180_ net98 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _0422_ _0531_ _2277_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4175_ _0784_ _0978_ _1089_ _0637_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3126_ _2421_ _2374_ _2423_ _2377_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3057_ _2271_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4263__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3369__A3 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _0967_ _0968_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3486__I _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3829__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4006__B2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3780__A3 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3517__B1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2740__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4955__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3296__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4931_ _1388_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ mod.registers.r6\[1\] _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3813_ _0651_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4548__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _1731_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2559__A1 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3744_ _0363_ _0372_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3220__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3675_ _0299_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2626_ _2006_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0232_ net78 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4720__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ mod.instr\[12\] _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5276_ _0163_ net99 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4227_ mod.ldr_hzd\[3\] _1235_ _1233_ mod.ldr_hzd\[1\] _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4484__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4158_ _0652_ _0706_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4089_ _0670_ _1085_ _1086_ _1098_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4711__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3278__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__I1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5336__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[4] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout110_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3460_ _0469_ _2327_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3075__B _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ _0393_ _0400_ _0401_ mod.registers.r1\[9\] _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ _0020_ net70 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__I _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _1868_ _1921_ _1922_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3269__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _0575_ _0642_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__A1 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2933__I _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A4 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4914_ _1313_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3441__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _1631_ _1749_ _1763_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _2385_ _1719_ _1721_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3727_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2952__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3658_ _2246_ _0661_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4796__S _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2609_ mod.pc_1\[4\] _1996_ _1994_ _1260_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3589_ _0550_ _0574_ _0589_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5328_ _0215_ net142 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _0146_ net90 mod.instr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4457__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4209__A1 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5359__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3432__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3983__A3 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2943__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3499__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2960_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__B1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2891_ _2187_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4630_ _1261_ _1575_ _1614_ _1599_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3187__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ _1525_ _1551_ _1553_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3584__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3512_ mod.registers.r7\[14\] _2169_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4492_ _2120_ _1391_ _1405_ _1384_ _1492_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_3443_ mod.registers.r2\[10\] _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ mod.pc_2\[9\] _2135_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5113_ _1923_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _1891_ _1898_ _1905_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_38_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3111__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3414__A2 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _1570_ _1749_ _1753_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3178__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ mod.registers.r3\[12\] _1707_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3193__A4 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4678__A1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2838__I _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_306 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4850__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3405__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4602__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2613__B1 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3341__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3090_ mod.registers.r7\[0\] _2168_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3644__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _2500_ _2529_ _0687_ _0355_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_62_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2943_ _2238_ _2188_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2874_ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4613_ _1265_ _1575_ _1598_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4544_ _1531_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4109__B1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3580__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1251_ _1477_ _1479_ _1321_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_89_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3426_ _0421_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout90_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__A3 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3332__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _2355_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3288_ _0284_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5027_ _1891_ _1892_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A1 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3399__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4060__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3946__I0 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3323__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__A1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3901__B _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_158 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_169 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4823__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2590_ _1987_ _1337_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3562__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ mod.pc_2\[2\] _1265_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4179__B _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3211_ _2382_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4191_ _1195_ _1200_ _1201_ _0652_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3865__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3142_ _2318_ _2435_ _2439_ mod.registers.r6\[1\] _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5067__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3073_ _2366_ _2368_ _2369_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_55_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3102__I mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3975_ _0626_ _0562_ _0840_ _0576_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4042__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2941__I mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2926_ _2221_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3258__B _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2857_ _2143_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2788_ _2100_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4527_ _1232_ _1519_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3772__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4458_ mod.pc_2\[13\] _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3305__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3409_ _0416_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4389_ mod.pc0\[10\] _1318_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5058__A1 _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2851__I _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4778__I _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3311__A4 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4024__A2 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _0698_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3783__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2586__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2711_ mod.des.des_dout\[8\] net4 _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3691_ _0699_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2642_ _1230_ _2015_ _2011_ mod.instr\[4\] _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3535__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4688__I _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _0248_ net147 mod.des.des_dout\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2573_ mod.des.des_dout\[16\] _1973_ _1974_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _0774_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5292_ _0179_ net102 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4243_ mod.pc_2\[6\] _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3838__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _0638_ _0947_ _1184_ _1164_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3125_ _2251_ _2375_ _2272_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5242__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3056_ _2313_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_36_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4263__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3958_ _0714_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2909_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3889_ _0326_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3526__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3829__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3451__B _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2782__S _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3214__B1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3765__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2568__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3517__B2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4190__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2740__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3296__A3 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2756__I _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3080__C _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4245__A2 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4930_ _1817_ _1818_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3587__I _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4861_ _1769_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3812_ _0822_ _0538_ _0815_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_20_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _1602_ mod.registers.r4\[7\] _1728_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2559__A2 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3743_ _0749_ _0750_ _0752_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3220__A3 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3674_ _2499_ _0680_ _0681_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ mod.pc_1\[11\] _2002_ _1932_ _1438_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4181__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ _0231_ net78 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2556_ _1967_ _1959_ _1968_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _0162_ net99 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ mod.instr_2\[5\] _1229_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4157_ _0463_ _0851_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3108_ _2191_ _2195_ _2198_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_83_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _1084_ _1097_ _0879_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3039_ _2322_ _2329_ _2336_ _2301_ mod.pc_2\[12\] _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__B1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3747__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3278__A3 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4475__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput14 io_in[5] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout103_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _2475_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ mod.pc\[13\] _1883_ _1884_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4011_ _2460_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3977__A1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4913_ _1793_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ mod.registers.r5\[11\] _1750_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3729__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _1540_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3726_ _0658_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2952__A2 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3657_ _2125_ _0639_ _0640_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4154__A1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2608_ _1812_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3588_ _0593_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3901__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _0214_ net142 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5258_ _0145_ net91 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ _2348_ _1216_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5189_ _0079_ net62 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4209__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3432__A3 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2640__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2943__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5303__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3408__B1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4454__C _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2890_ _2124_ _2127_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2631__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2919__C1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ mod.registers.r1\[1\] _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3187__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ mod.registers.r1\[14\] _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4491_ _1412_ _2346_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4136__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3442_ mod.registers.r4\[10\] _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3814__B _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3373_ _0379_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ mod.instr\[9\] _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1902_ _1907_ _1841_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3105__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3111__A2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__B _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3414__A3 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4611__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ mod.registers.r5\[4\] _1750_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3178__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _1632_ _1706_ _1708_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3709_ _0716_ _0718_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4689_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4127__A1 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3724__B _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_307 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4850__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2861__A1 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2861__B2 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4989__I0 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__A1 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__B2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4366__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4669__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _1000_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2942_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2873_ _2152_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _1531_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ mod.pc_2\[0\] _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4109__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3580__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _1251_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3425_ _0422_ _2245_ _2247_ _2241_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__3332__A2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3356_ _0366_ _0310_ _0314_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout83_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3287_ _0294_ _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _1891_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4832__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3399__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4596__A1 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__A3 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3946__I1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3323__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4520__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3874__A3 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_159 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__B1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3210_ mod.registers.r3\[3\] _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4511__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ _0820_ _0742_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3141_ _2174_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2695__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3072_ _2193_ _2362_ _2214_ mod.registers.r1\[0\] _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_55_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3078__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4195__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3974_ _0836_ _0837_ _0576_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2925_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2856_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5171__CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2787_ net3 mod.des.des_dout\[23\] _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4526_ mod.rd_3\[0\] _1513_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4457_ _1460_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3305__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3408_ _0417_ _2509_ _2317_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_58_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4388_ mod.pc\[10\] _1351_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ _0333_ _0337_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4805__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ _1876_ _1878_ _1319_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3241__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3792__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4741__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5049__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3203__I mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2807__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3480__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4024__A3 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5194__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3078__C _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout133_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _2043_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3783__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3690_ _0408_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4969__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2641_ _1796_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3535__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2572_ mod.instr\[16\] _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5360_ _0247_ net143 mod.des.des_dout\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4311_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ _0178_ net101 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4242_ _2349_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3299__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__B _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4173_ _1056_ _0923_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3124_ _2195_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout46_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3471__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__B _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ _0501_ _0507_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2908_ mod.instr_2\[12\] _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4971__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3888_ _0604_ _0692_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2982__B1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2839_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _1423_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3023__I mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3462__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2862__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__A1 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3693__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4714__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3517__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4190__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3296__A4 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3453__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3868__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4860_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3811_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3205__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _0272_ _1719_ _1730_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3742_ _0634_ _0622_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3673_ _0683_ _2527_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4705__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2624_ _2005_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _0230_ net62 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4181__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2555_ mod.des.des_dout\[11\] _1962_ _1963_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _0161_ net121 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__I _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4225_ mod.ldr_hzd\[4\] _1231_ _1233_ mod.ldr_hzd\[5\] mod.ldr_hzd\[7\] _1235_ _1236_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4156_ _0992_ _0865_ _0978_ _0835_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_68_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3692__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3107_ mod.registers.r2\[1\] _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4087_ _1084_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3038_ _2135_ _2333_ _2334_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4989_ _1387_ _1393_ _1209_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4172__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3278__A4 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3683__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2793__S _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput15 io_in[6] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4312__I _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4010_ _0616_ _0744_ _0677_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3674__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3426__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4912_ _1226_ _1799_ _1804_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__A2 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4843_ _0438_ _1746_ _1762_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__A2 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _1717_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3725_ _0547_ _0667_ _0672_ _0735_ _0721_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3656_ _0600_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4154__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2607_ _1995_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3587_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5326_ _0213_ net84 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3901__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _0144_ net91 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4208_ _1216_ mod.ldr_hzd\[4\] _2348_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3665__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5188_ _0078_ net62 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _0575_ _0885_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3301__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5255__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2928__B1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3423__A4 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2919__B1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2919__C2 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3187__A3 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3510_ _0519_ _2509_ _2327_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4490_ _1491_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4136__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3441_ _0451_ _2509_ _2320_ _0438_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3372_ _2300_ _0380_ _0381_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5111_ _1958_ _1959_ _1960_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _1865_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5128__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3111__A3 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4072__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4661__B _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2960__I _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4826_ _1565_ _1749_ _1752_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3178__A3 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ mod.registers.r3\[11\] _1707_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3708_ _0537_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4688_ _1662_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__I _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3639_ _0648_ _2261_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_122_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3886__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__A2 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5309_ _0196_ net88 mod.instr_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_308 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4686__I0 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4989__I1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3810__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2870__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4366__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3915__B _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A1 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4465__C _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3990_ _0351_ _0907_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2941_ mod.instr_2\[1\] _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3801__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4481__B _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2872_ mod.registers.r7\[15\] _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _1586_ _1284_ _1587_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _2130_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4473_ _1416_ _0932_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3424_ _0368_ _0427_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3355_ _0364_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3332__A3 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout76_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3286_ _2542_ _2453_ _0296_ _2445_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2955__I _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ mod.pc\[8\] _1346_ _1334_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4596__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4809_ _0525_ _1719_ _1740_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3323__A3 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4520__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3026__I _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2865__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__A1 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__A2 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4036__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4339__A2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3140_ mod.registers.r7\[1\] _2437_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ _2367_ _2196_ _2357_ mod.registers.r6\[0\] _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3078__A2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4195__C _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _0825_ _0827_ _0601_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _2194_ _2206_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3250__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2855_ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5316__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2786_ _2089_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4525_ _1511_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2761__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4456_ _1143_ _1156_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3407_ mod.registers.r1\[11\] _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4502__A2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4387_ mod.pc0\[3\] _1249_ _1389_ _1348_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _2461_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3269_ _2493_ _2152_ _2175_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4266__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5008_ _1863_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4405__I _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3241__A2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4741__A2 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__S _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2595__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3359__C _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2640_ _1989_ _2014_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout126_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3535__A3 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ _1978_ _1970_ _1979_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4310_ _1208_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3940__B1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5290_ _0177_ net101 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ mod.pc_2\[7\] _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3299__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4172_ _1176_ _1178_ _0822_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3123_ mod.instr_2\[4\] _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4248__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3054_ _2338_ _2351_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4934__B _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout39_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3956_ _0754_ _0755_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4420__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3223__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2907_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3887_ _0642_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2982__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2838_ _2135_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2982__B2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4723__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2769_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4508_ _1460_ _1197_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _1398_ _1442_ _1444_ _1288_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4239__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3462__A2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3214__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4411__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__A2 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4175__B1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4714__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3773__I0 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4478__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5161__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3453__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _0820_ _0653_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4790_ _1593_ _1720_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4402__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3205__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3741_ _0751_ _0686_ _0328_ _0687_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3672_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ mod.pc_1\[10\] _2002_ _2000_ _1399_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4705__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5342_ _0229_ net147 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2554_ mod.instr\[11\] _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4929__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5273_ _0160_ net122 mod.pc0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _0844_ _0805_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3106_ _2355_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4086_ _1065_ _0903_ _0905_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2963__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3037_ _2288_ _2290_ _2296_ mod.registers.r4\[12\] _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3444__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2652__B1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4988_ _1854_ _1860_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3939_ _0606_ _0567_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3380__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3132__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5184__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3034__I _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2873__I _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3199__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 io_in[7] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4699__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3879__I _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3426__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4623__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4911_ mod.rd_3\[1\] _1800_ _1802_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ _1623_ _1743_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3729__A3 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4926__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ _0722_ _0731_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _0628_ _0633_ _0644_ _0647_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_2606_ mod.pc_1\[3\] _1990_ _1994_ mod.pc_2\[3\] _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3586_ _0594_ _0595_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3362__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2958__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ _0212_ net84 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4378__C _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5256_ _0143_ net111 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4207_ _0422_ mod.ldr_hzd\[5\] _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5187_ _0077_ net39 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3665__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ _0874_ _1148_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ _0902_ _0801_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4614__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2625__B1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__A3 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4090__A2 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__B1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2928__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2928__B2 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3353__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2868__I mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4853__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3408__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2616__B1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2552__B _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2919__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2919__B2 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3187__A4 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3440_ mod.registers.r3\[10\] _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3344__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3371_ _2180_ _0375_ _2519_ mod.registers.r4\[9\] _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_124_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3895__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5110_ mod.des.des_dout\[8\] _1951_ _1952_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _1899_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4844__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4942__B _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ mod.registers.r5\[3\] _1750_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5021__A1 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3178__A4 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _1688_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3707_ _2311_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _1664_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3638_ _0595_ mod.funct3\[0\] _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3335__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3569_ _2137_ _2185_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5064__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _0195_ net104 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__A1 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5239_ _0126_ net124 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_309 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4835__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3638__A2 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4686__I1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2697__I0 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5222__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3271__B1 _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5372__CLK net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4118__A3 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2598__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3877__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A2 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4318__I _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ mod.funct7\[2\] _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2871_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4610_ _1252_ _1544_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4541_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4472_ _1254_ _1255_ _1279_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__3317__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3423_ _0430_ _0431_ _0432_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4002__B _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3354_ mod.pc_2\[5\] _2301_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ mod.funct3\[1\] _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5245__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout69_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__A2 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2971__I _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4808_ _1651_ _1720_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3556__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4898__I _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _1566_ _1693_ _1697_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3323__A4 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3751__B _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4808__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4284__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3926__B _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3217__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5268__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__C _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3070_ _2367_ _2213_ _2208_ mod.registers.r5\[0\] _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _0578_ _0871_ _0982_ _0882_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2923_ _2192_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2854_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2785_ _2098_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4455_ _1416_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ mod.registers.r3\[11\] _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4386_ _1348_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2966__I _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ mod.funct7\[1\] _2240_ _2339_ _2404_ _0342_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_4
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3268_ mod.registers.r3\[6\] _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__S _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4266__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _1870_ _1875_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3199_ _2134_ _2491_ _2492_ _2496_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3777__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5010__C _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3241__A3 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3701__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4257__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3465__B1 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ mod.des.des_dout\[15\] _1973_ _1974_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3940__B2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3299__A3 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2786__I _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4171_ _0743_ _1181_ _0734_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3122_ _2414_ _2416_ _2417_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_68_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4248__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__S _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3053_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3471__A3 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3759__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3955_ _0759_ _0502_ _0936_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4950__B _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4420__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3223__A3 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ mod.instr_2\[13\] _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3886_ _0686_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2982__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2837_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4241__I mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2768_ mod.des.des_counter\[2\] _1411_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4507_ _2120_ _1499_ _1501_ _1195_ _1503_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_2699_ mod.des.des_dout\[3\] net16 _2044_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4438_ _1398_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4487__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4369_ _1373_ _1374_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3462__A3 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4416__I _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2670__A1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2973__A2 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4175__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3773__I1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4478__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5306__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2555__B _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A1 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__B2 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4402__A2 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _0357_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3671_ _2258_ _2481_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2622_ _2004_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3913__A1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2553_ _1965_ _1959_ _1966_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5341_ _0228_ net148 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4181__A4 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5272_ _0159_ net121 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4469__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ mod.instr_2\[4\] mod.instr_2\[3\] _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4154_ _0959_ _1117_ _0953_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3105_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4085_ _1084_ _0802_ _0803_ _0625_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3036_ _2331_ mod.registers.r3\[12\] _2146_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2652__B2 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ mod.pc\[2\] _1844_ _1857_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3938_ _0576_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3869_ _0790_ _0878_ _0879_ _0795_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_109_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4157__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3904__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3743__C _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5329__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5016__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3132__A2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2891__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3435__A3 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3050__I _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2643__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4590__B _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 io_in[8] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4148__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3225__I mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4320__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4871__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__B1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4623__A2 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ _1232_ _1799_ _1803_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _0387_ _1746_ _1761_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4387__A1 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4387__B2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4772_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3723_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4139__A1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3654_ _0543_ _0651_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2605_ _1931_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3585_ mod.funct3\[0\] _2260_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3362__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5324_ _0211_ net84 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout99_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _0142_ net109 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3114__A2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ mod.ldr_hzd\[0\] mod.ldr_hzd\[1\] mod.ldr_hzd\[2\] mod.ldr_hzd\[3\] _1216_
+ _0428_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5186_ _0076_ net80 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3665__A3 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2974__I _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _0808_ _0950_ _1144_ _1145_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_96_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _0338_ _0349_ _0891_ _0657_ _0848_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4614__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__B2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__B2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2928__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4066__B1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2616__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2616__B2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2919__A2 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4479__C _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout101_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3344__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3370_ _2149_ mod.registers.r3\[9\] _2146_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5040_ _1407_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3280__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4514__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _1559_ _1749_ _1751_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5021__A2 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _1689_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3706_ _2312_ _0585_ _2351_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4780__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _1660_ mod.registers.r2\[0\] _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2969__I _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3637_ _0594_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3293__C _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3335__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3568_ _2379_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _0194_ net110 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3499_ _2338_ _2350_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3099__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _0125_ net123 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4835__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2846__A1 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _0059_ net51 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2697__I1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__A3 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5012__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2879__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3014__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _1531_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4762__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ mod.pc0\[6\] _1309_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3317__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3422_ _0393_ _0400_ _0401_ mod.registers.r1\[11\] _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3353_ _0319_ _0323_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3614__S _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3284_ _2256_ _2271_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _1862_ _1877_ _1881_ _1887_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3253__A1 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ _1646_ _1735_ _1739_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2999_ _2288_ _2172_ _2296_ mod.registers.r6\[13\] _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4753__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ mod.registers.r3\[3\] _1694_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _1536_ _1502_ _1576_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3483__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _0583_ _0861_ _0863_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3235__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2922_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2853_ mod.instr_2\[10\] _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4735__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2784_ net2 mod.des.des_dout\[22\] _2094_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _1226_ _1513_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4454_ _1317_ _1449_ _1458_ _1356_ _1459_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4948__B _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3405_ _0415_ _2510_ _2483_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4385_ _1283_ _1390_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout81_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3336_ _0343_ _0344_ _0345_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_112_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3267_ _0274_ _0275_ _0276_ _0277_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5006_ _1850_ _1874_ _1870_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3198_ _2494_ _2326_ _2495_ mod.registers.r2\[2\] _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3299__B _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3226__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3241__A4 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__I _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3762__B _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3162__B1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3053__I _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3465__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3465__B2 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3480__A4 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4612__I _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4170_ _0751_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3121_ _2408_ _2415_ _2418_ mod.registers.r1\[1\] _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_95_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3052_ _2342_ _2347_ _2349_ _2309_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3471__A4 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4956__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ _0944_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3223__A4 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3847__B _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2905_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3885_ _0890_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2836_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2767_ _1657_ _2081_ _2087_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4506_ _1423_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2698_ _2047_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _0976_ _0999_ _1322_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4368_ _1327_ _1328_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3319_ _2428_ _2484_ _2392_ mod.registers.r1\[4\] _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ mod.pc0\[0\] _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3447__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4633__S _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4947__A1 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5258__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4175__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__I1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3686__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3989__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4938__A1 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3670_ _0673_ _0354_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4166__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2621_ mod.pc_1\[9\] _2002_ _2000_ _1373_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5340_ _0227_ net147 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2552_ mod.des.des_dout\[10\] _1962_ _1963_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5271_ _0158_ net111 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ mod.instr_2\[4\] _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2724__I0 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4153_ _0790_ _0921_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3104_ _2386_ _2389_ _2399_ _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _0675_ _0849_ _0852_ _0904_ _0732_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_110_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3035_ _2331_ _2332_ _2296_ mod.registers.r2\[12\] _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_290 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout44_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _1309_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3937_ _0785_ _0618_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3601__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3868_ _0669_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4157__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2819_ _2118_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3799_ _0632_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5106__A1 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5083__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2715__I0 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3132__A3 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2891__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3435__A4 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__A2 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 io_in[9] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4148__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__A3 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4337__I _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__B2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4840_ _1616_ _1757_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4387__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4771_ _1713_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3722_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4005__C _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3653_ _0542_ _0656_ _0659_ _0660_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4800__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2604_ _1993_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3584_ mod.funct3\[1\] _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5323_ _0210_ net81 mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2570__A1 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5254_ _0141_ net112 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ _0401_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5185_ _0075_ net80 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4136_ _0550_ _0946_ _1146_ _0631_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _1073_ _1077_ _0776_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3018_ _2140_ _2315_ _2155_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2990__I _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _1318_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5078__I _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout151 net1 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3510__B1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3061__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4066__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__B2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3010__B _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2552__A1 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3280__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4823_ mod.registers.r5\[2\] _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5319__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _0451_ _1690_ _1705_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3705_ _0703_ _0713_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3855__B _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__A2 _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4530__I _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3636_ _0541_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3567_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3146__I mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5306_ _0193_ net109 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3498_ _2338_ _2350_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5237_ _0124_ net128 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3099__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5168_ _0058_ net57 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4119_ _1065_ _0903_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4048__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _1801_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__S _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4220__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__I _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4615__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3798__B1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3014__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4350__I _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4470_ mod.pc\[6\] _1351_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ _0423_ _0400_ _0401_ mod.registers.r5\[11\] _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3352_ _0357_ _0358_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3283_ _2377_ _0288_ _0293_ _2341_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_98_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5022_ _1865_ _1888_ _1889_ _1847_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5141__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3789__B1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3253__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4450__A1 mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ mod.registers.r4\[13\] _1736_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3005__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4737_ _1560_ _1693_ _1696_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4753__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4668_ mod.des.des_dout\[32\] _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3619_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4505__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4599_ _1532_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4269__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3180__A1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3483__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ _0979_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3235__A2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2921_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2852_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4735__A2 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2783_ _2097_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4522_ mod.rd_3\[1\] _1513_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4453_ _2534_ _2540_ _1385_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3404_ mod.registers.r4\[11\] _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4384_ _1359_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3335_ mod.registers.r7\[4\] _2365_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3266_ _2148_ _2546_ _2155_ mod.registers.r1\[6\] _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5005_ _1873_ _1454_ _1209_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3197_ _2395_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3226__A2 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4423__A1 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2704__S _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2737__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3934__B1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5187__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__B _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4111__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3465__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4662__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2673__B1 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4178__B1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3509__I mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2728__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3244__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _2207_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3051_ _2348_ _2275_ _2276_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4653__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ _2264_ _0939_ _0945_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2904_ mod.instr_2\[14\] _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3884_ _0893_ _0894_ _0328_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _2131_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2766_ mod.registers.r7\[15\] _2082_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4505_ _1460_ _0889_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2697_ mod.des.des_dout\[2\] net15 _2044_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _1437_ mod.pc_2\[12\] _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _1375_ _1331_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4892__A1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3318_ _2494_ _2394_ _2495_ mod.registers.r2\[4\] _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_59_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _1248_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3249_ _2148_ _2546_ _2441_ mod.registers.r1\[7\] _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_58_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3447__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4644__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2655__B1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3329__I mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__A1 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3064__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3686__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4635__A1 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4938__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__A1 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3997__I0 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5352__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2620_ _2003_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3374__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ mod.instr\[10\] _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ _0157_ net111 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5115__A2 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3126__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _2372_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3677__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2724__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4152_ _0743_ _1162_ _0734_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3103_ _2400_ _2265_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4083_ _1088_ _1093_ _0777_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3034_ _2326_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2637__B1 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_280 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_291 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__B _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout37_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4929__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _1850_ _1856_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5051__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _0592_ _0806_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2818_ _2116_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3798_ _0625_ _0805_ _0808_ _0613_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3365__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2988__I mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2749_ _2065_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3380__A4 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4419_ _1416_ _0813_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_120_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4865__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2715__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A2 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3059__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4111__C _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3371__A4 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3108__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2706__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2619__B1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4770_ _1518_ _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ _0648_ _2254_ _0657_ _2261_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2802__S _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3652_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2603_ mod.pc_1\[2\] _1990_ _1933_ _1264_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3583_ mod.funct3\[2\] _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3898__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ _0209_ net82 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _0140_ net113 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4847__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5248__CLK net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4204_ _2126_ _1213_ _1214_ _2181_ _2247_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_87_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5184_ _0074_ net80 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4135_ _0627_ _0948_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__I _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ _0947_ _0995_ _1076_ _0635_ _0924_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4075__A2 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3017_ _2160_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _1369_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _0599_ _0846_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4899_ _1795_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3338__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__I _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout130 net131 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout141 net151 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__B _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3510__B2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4066__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3010__C _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3577__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2552__A2 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3501__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__A2 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3280__A3 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _1745_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4753_ _1623_ _1691_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _2313_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4684_ _1515_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__B _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3635_ _2253_ _0645_ _0596_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_127_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5305_ _0192_ net90 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3497_ _0501_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5236_ _0123_ net126 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3099__A3 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _0057_ net54 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4118_ _2263_ _0749_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5098_ _1924_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input17_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4049_ _1054_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__B _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3420_ _0397_ _0428_ _0429_ mod.registers.r6\[11\] _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3351_ _0361_ _2541_ _2544_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3282_ _0289_ _0290_ _0291_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ mod.pc\[7\] _1866_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3710__I _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ _1639_ _1735_ _1738_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2997_ _2174_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4736_ mod.registers.r3\[2\] _1694_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3157__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _1552_ _1646_ _1647_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3618_ _2507_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4598_ _1527_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3713__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3549_ _2404_ _0311_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4269__A2 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _0106_ net103 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3952__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3067__I _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3180__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3530__I _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2691__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3235__A3 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2920_ _2202_ _2194_ _2206_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_31_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2851_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4361__I _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2782_ net18 mod.des.des_dout\[21\] _2094_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3943__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4521_ _1507_ _1512_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ mod.pc0\[5\] _1369_ _1455_ _1338_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__I0 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _0410_ _0411_ _0412_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4383_ _1172_ _1101_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _2361_ _2362_ _2357_ mod.registers.r4\[4\] _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3265_ mod.registers.r7\[6\] _2437_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4120__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5004_ _1856_ _1861_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3196_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout67_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4671__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2809__I0 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2985__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4204__C _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1639_ _1670_ _1684_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2720__S _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3615__I _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2673__A1 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2673__B2 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4178__A1 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__B2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__C _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5131__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3525__I _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3050_ _2205_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4356__I _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _0933_ _0651_ _0952_ _0632_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2903_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3883_ _0609_ _0349_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2834_ mod.instr_2\[2\] mod.instr_2\[0\] _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3916__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2765_ _2086_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1213_ _2117_ _1205_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2696_ _2046_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4435_ _1436_ _1438_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3144__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4366_ mod.pc_2\[8\] _1328_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3317_ _0326_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _1301_ _1305_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3248_ _2160_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3447__A3 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4644__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3170__I mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2655__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3179_ _2473_ mod.registers.r3\[2\] _2222_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_66_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2655__B2 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2715__S _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3080__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5154__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__A1 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__I0 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3135__A2 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4635__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2646__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__B1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3997__I1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__B _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3374__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4323__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4220_ _1230_ mod.instr_2\[3\] _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _0465_ _0769_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2885__A1 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3102_ mod.pc_2\[0\] _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _0977_ _1089_ _1090_ _1091_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3033_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2637__A1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_270 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2637__B2 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_281 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_292 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _1850_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3935_ _0611_ _0624_ _0843_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3062__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5177__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3866_ _0683_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2817_ mod.des.des_counter\[1\] _0000_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3797_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3365__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2748_ _2076_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2679_ _2037_ _2038_ _1815_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4418_ mod.pc\[11\] _1348_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _1264_ _1265_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_113_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A3 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4305__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3803__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2867__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__B2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3292__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _0544_ _0535_ _0730_ _0671_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _2252_ _0649_ _2268_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2602_ _1992_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3582_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ _0208_ net81 mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5252_ _0139_ net101 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4847__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ mod.ldr_hzd\[0\] mod.ldr_hzd\[1\] mod.ldr_hzd\[2\] mod.ldr_hzd\[3\] _2164_
+ _2154_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5183_ _0073_ net77 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _0584_ _0587_ _0992_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4065_ _1074_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3869__B _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3016_ mod.registers.r1\[12\] _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3283__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4544__I _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4967_ mod.pc\[0\] _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3918_ _0686_ _0651_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4783__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4898_ _1795_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3849_ _0603_ _0858_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3338__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4838__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout120 net125 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3623__I _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout142 net144 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3510__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3265__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2593__B _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4364__I mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3280__A4 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4821_ _1745_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4752_ _1704_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4765__A1 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3703_ _0511_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _1518_ _1521_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3634_ _2254_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5215__CLK net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3565_ _0551_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _0191_ net90 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout97_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3496_ _0502_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5365__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5235_ _0122_ net118 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3099__A4 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _0056_ net43 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4117_ _2460_ _2463_ _2499_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ mod.instr\[5\] _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _1055_ _1058_ _0598_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3256__A1 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5310__D _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3008__A1 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3008__B2 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3618__I _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4508__A1 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3731__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4449__I _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3495__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A3 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3183__B1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3350_ _0359_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _2367_ _2196_ _2357_ mod.registers.r6\[6\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _1886_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3789__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4986__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3253__A4 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4738__A1 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4804_ mod.registers.r4\[12\] _1736_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4822__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2996_ _2288_ _2290_ _2293_ mod.registers.r5\[13\] _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3005__A4 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _1551_ _1693_ _1695_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__B _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3410__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4666_ mod.registers.r1\[13\] _1526_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4978__B _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3617_ _0613_ _0625_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4597_ _1531_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3713__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4910__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3548_ _0557_ _0558_ _2131_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _0477_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5218_ _0105_ net103 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3477__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ _0039_ net72 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__I _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3401__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__C _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3083__I mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3180__A3 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5215__D _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4907__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3811__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3235__A4 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2850_ _2139_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout147_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2781_ _2096_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _2375_ _1500_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3943__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4451_ _1364_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ _2331_ _2332_ _2296_ mod.registers.r2\[11\] _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4743__I1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4382_ _2523_ _1262_ _1273_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_98_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2754__I0 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ _2193_ _2213_ _2208_ mod.registers.r1\[4\] _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ _2179_ _2152_ _2439_ mod.registers.r6\[6\] _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3459__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ mod.pc\[5\] _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3195_ _2138_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2682__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__A1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2809__I1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A3 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4552__I _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2979_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3934__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4718_ mod.registers.r2\[12\] _1671_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4649_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3698__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2745__I0 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__I _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3631__I _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3870__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2673__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4178__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3925__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2728__A3 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2710__I _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3541__I _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3861__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3208__A4 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3697__B _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3951_ _0795_ _0960_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2902_ _2193_ _2196_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_31_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ _0748_ _0750_ _0892_ _0753_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4169__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2833_ mod.instr_2\[1\] _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ _1652_ mod.registers.r7\[14\] _2077_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4503_ _1207_ _1312_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3716__I _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2695_ mod.des.des_dout\[1\] net14 _2044_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2620__I _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4434_ _1439_ _1429_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4365_ _0532_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3316_ _0324_ _0310_ _0314_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1300_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3247_ mod.registers.r7\[7\] _2437_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3447__A4 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3178_ _2473_ _2474_ _2475_ mod.registers.r1\[2\] _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_67_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__S _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3626__I _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__I1 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3135__A3 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4332__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3843__B2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3071__A2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4571__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4150_ _1159_ _1160_ _0671_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3101_ _2390_ _2393_ _2397_ _2398_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ _0792_ _1034_ _0920_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4087__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3032_ _2139_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_260 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2637__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_271 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_282 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_293 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _1855_ _1362_ _1320_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3934_ _0709_ _0850_ _0853_ _0707_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3062__A2 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3865_ _0857_ _0865_ _0873_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4830__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ _2113_ mod.des.des_counter\[0\] _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _0593_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ _1601_ mod.registers.r7\[7\] _2066_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3365__A3 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2678_ mod.valid_out3 _1814_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4417_ _1350_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4348_ _1267_ _1269_ _1270_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4277__I _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4279_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2726__S _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5121__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4002__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5271__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2564__A1 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3108__A3 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4305__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3816__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2619__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3292__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4616__I0 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3650_ _2256_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ mod.pc_1\[1\] _1990_ _1933_ mod.pc_2\[1\] _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3581_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ net311 net81 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _0138_ net113 mod.valid1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3504__B1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4202_ _2187_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _0072_ net39 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4133_ _0555_ _0572_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4064_ _0553_ _0825_ _0833_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _2311_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3283__A2 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__I0 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5294__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3035__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4232__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4966_ _1472_ _1840_ _1841_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3917_ _0737_ _0693_ _0927_ _0851_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4783__A2 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4897_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _0831_ _0832_ _0268_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_20_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3779_ _2159_ _2165_ _2170_ _2184_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_164_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout110 net112 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2849__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout132 net133 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__C _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5167__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3265__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ _1550_ _1746_ _1748_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__B2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4751_ _1617_ mod.registers.r3\[9\] _1699_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4380__I _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2776__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ _0705_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ _1540_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _0637_ _0638_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3564_ _0563_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _0190_ net84 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3495_ _0408_ _0504_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _0121_ net117 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _0055_ net72 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4116_ _0844_ _0803_ _1126_ _0662_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5096_ _1947_ _1948_ _1949_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4047_ _0805_ _1057_ _0981_ _0882_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_44_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3008__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4949_ mod.pc_1\[7\] _1827_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4290__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2767__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3495__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4692__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3247__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__A2 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2758__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3972__C _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3183__A1 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3183__B2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2930__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3280_ _2269_ _2422_ _2536_ mod.registers.r2\[6\] _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4375__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _1632_ _1735_ _1737_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4738__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2995_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4734_ mod.registers.r3\[1\] _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3410__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4665_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5332__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3882__C _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3616_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4596_ mod.des.des_dout\[24\] _1542_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3547_ _2366_ _2368_ _2369_ _2370_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4910__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3478_ _0486_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5217_ _0104_ net113 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3477__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _0038_ net70 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4285__I _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _1936_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3401__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3165__A1 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3180__A4 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3468__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5205__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5355__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2780_ net17 mod.des.des_dout\[20\] _2094_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4450_ mod.pc\[5\] _1365_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3156__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3401_ _2517_ _2290_ _2293_ mod.registers.r5\[11\] _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4381_ _1387_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2754__I1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3332_ _2221_ mod.registers.r3\[4\] _2359_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_112_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ _2179_ _2546_ _2441_ mod.registers.r5\[6\] _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3459__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4200__S0 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4656__A1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5002_ _1868_ _1871_ _1872_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3194_ _2488_ _2326_ _2295_ mod.registers.r6\[2\] _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4833__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2978_ _2238_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3395__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _1632_ _1670_ _1683_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ mod.des.des_dout\[29\] _1626_ _1628_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _0607_ _1529_ _1546_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3698__A2 _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2745__I1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2658__B1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5072__A1 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3138__A1 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__A1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3310__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _0776_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2901_ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3881_ _0609_ _0793_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4574__B1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2763_ _1645_ _2081_ _2085_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2901__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4502_ _2364_ _2371_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2694_ _2045_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3129__A1 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _1436_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3144__A4 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4364_ mod.pc_2\[9\] _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3315_ _0310_ _0314_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_98_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3732__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4295_ _2400_ _1266_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3246_ _2542_ _2464_ _2543_ _2445_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA_fanout72_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ _2207_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5054__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4563__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4868__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3135__A4 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3540__A1 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A1 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3089__I mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3071__A3 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3359__A1 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3359__B2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4020__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3980__C _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3552__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ _2141_ _2171_ _2396_ mod.registers.r2\[0\] _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2885__A3 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _0949_ _1031_ _0881_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3031_ _2323_ _2327_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_250 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_261 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_272 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_283 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_294 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3501__B _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3047__B1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ mod.pc\[2\] _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3598__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3933_ _0814_ _0939_ _0941_ _0943_ _0772_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_51_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3062__A3 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3864_ _0629_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2815_ _2115_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _0548_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3727__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2746_ _2075_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3365__A4 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3770__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2677_ mod.valid2 _1823_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4416_ _2116_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3522__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4558__I _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4347_ _2119_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3229_ _2498_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2867__A3 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4069__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4616__I1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4136__C _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4931__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4152__B _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout122_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _1991_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3580_ mod.funct7\[0\] _0368_ _0590_ _2245_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3752__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2555__A2 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _0137_ net127 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3504__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4201_ _2150_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _0071_ net68 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4132_ _0767_ _1139_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4063_ _0602_ _0830_ _0859_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3014_ _2307_ _2310_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4327__B _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3283__A3 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__I1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _1805_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3035__A3 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3916_ _0691_ _0692_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4896_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3847_ _0789_ _0829_ _0476_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_164_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ _0608_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3743__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2729_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout100 net101 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout111 net112 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout122 net124 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout133 net134 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3125__C _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout144 net150 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3982__A1 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4198__I _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4147__B _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ _1703_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3701_ _0704_ _0499_ _0706_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3973__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _1552_ _1658_ _1659_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3632_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3563_ _0555_ _0567_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5302_ _0189_ net105 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3494_ _0386_ _0404_ _0406_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_103_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _0120_ net117 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5164_ _0054_ net58 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ _1065_ _0650_ _1124_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ mod.des.des_dout\[4\] _1940_ _1941_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5261__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ _0840_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4453__A2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _1475_ _1830_ _1829_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4879_ _1609_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5005__I1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4141__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4692__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3650__I _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5134__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3183__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__S _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2930__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4683__A2 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__I mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2904__I mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ mod.registers.r4\[11\] _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2994_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4733_ _1688_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4664_ mod.des.des_dout\[31\] _1626_ _1642_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3615_ _2482_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4595_ _1583_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3174__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4371__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3546_ _2358_ _2360_ _2363_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ _2455_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4123__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _0002_ _0006_ net146 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_88_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4674__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5147_ _0037_ net70 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2685__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _1923_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input15_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4426__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _0356_ _0373_ _0936_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_37_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5157__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2750__S _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3401__A3 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3645__I _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3165__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4362__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2676__A1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3476__I0 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__B1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__B _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3156__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ _2180_ _2153_ _2519_ mod.registers.r6\[11\] _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4353__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4380_ _1313_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ _0339_ _2467_ _2406_ _0340_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_98_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3262_ _0272_ _2384_ _2299_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4200__S1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4656__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ mod.pc\[4\] _1865_ _1802_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3290__I _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3193_ _2488_ _2484_ _2392_ mod.registers.r5\[2\] _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320__311 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4408__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2634__I _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3919__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2977_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3395__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ mod.registers.r2\[11\] _1671_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4070__B _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4647_ _1535_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4578_ _1547_ _1493_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3698__A3 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3529_ _2185_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4647__A2 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2658__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2658__B2 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2745__S _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5072__A2 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3138__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4335__A1 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2719__I _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2649__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3310__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2900_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _0608_ _0350_ _0348_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3994__B _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _2126_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4574__A1 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__B2 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2762_ mod.registers.r7\[13\] _2082_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _0001_ _1478_ _1498_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2693_ mod.des.des_dout\[0\] net13 _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3129__A2 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4326__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ mod.pc_2\[11\] _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4363_ _1370_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2888__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3314_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _1302_ _1115_ _1304_ _0740_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4629__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3245_ _2251_ _2273_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3176_ _2204_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3065__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4565__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4868__A2 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5045__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3056__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3071__A4 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3359__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3531__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2885__A4 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3030_ mod.registers.r7\[12\] _2169_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xtiny_user_project_240 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3295__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_251 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4492__B1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_262 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_273 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_284 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_295 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3501__C _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3047__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3047__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ _0759_ _0942_ _0898_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3863_ _0594_ _0595_ _0596_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_31_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__I _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2814_ net130 _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5218__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3794_ _0629_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2745_ _1594_ mod.registers.r7\[6\] _2066_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3944__S _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3770__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ _2032_ _2036_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4415_ mod.pc0\[4\] _1369_ _1419_ _1338_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5368__CLK net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3522__A2 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4346_ _1317_ _1337_ _1354_ _0001_ _1355_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_87_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _1210_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3899__B _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ _2507_ _2525_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3159_ _2300_ _2436_ _2440_ _2442_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3038__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4710__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3513__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2867__A4 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3277__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3292__A4 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3029__A1 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4529__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3201__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout115_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ mod.ldr_hzd\[4\] mod.ldr_hzd\[5\] mod.ldr_hzd\[6\] mod.ldr_hzd\[7\] _2164_
+ _2154_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3504__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _0070_ net58 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _0767_ _1141_ _0734_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _0807_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3013_ _2307_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3939__S _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4964_ mod.pc_1\[13\] _1806_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3035__A4 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _0915_ _0925_ _0778_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4895_ _1507_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3846_ _0804_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ _0631_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2728_ _1517_ _1522_ _1715_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2659_ _2025_ _2026_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout101 net102 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout112 net115 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4329_ _1302_ _1039_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout134 mod.clk net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout145 net149 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3259__A1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4759__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2793__I0 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3383__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3498__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3558__I _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _0463_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3973__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4680_ mod.registers.r1\[15\] _1526_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3725__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3562_ _0555_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5301_ _0188_ net109 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2784__I0 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3493_ _0503_ _0486_ _0488_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5232_ _0119_ net119 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3489__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5163_ _0053_ net73 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4114_ _0804_ _0619_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5094_ _1936_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4045_ _0569_ _0843_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ mod.pc_1\[6\] _1827_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3413__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4878_ _1769_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ _2400_ _0789_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4429__B1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3378__I _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3183__A3 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4937__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3643__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4672__I _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4801_ _1717_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2993_ _2143_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4732_ _1689_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4663_ _1535_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3614_ _0618_ _0624_ _0577_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4594_ _1581_ mod.registers.r1\[5\] _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3545_ mod.pc_2\[9\] _2136_ _0379_ _0383_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3476_ mod.funct7\[0\] _2293_ _2274_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5215_ _0001_ _0005_ net146 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__4123__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5146_ _0036_ net67 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2685__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ mod.instr\[0\] _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4028_ _0818_ _1024_ _1029_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3937__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3401__A4 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4362__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3476__I1 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__C _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4050__B2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5251__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _2203_ _2422_ _2536_ mod.registers.r6\[4\] _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3261_ mod.registers.r4\[6\] _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3571__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3313__B1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5000_ _1863_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3192_ _2485_ _2486_ _2487_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3864__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2915__I _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3947__S _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2976_ _2273_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _0454_ _1666_ _1682_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3746__I _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4646_ _1255_ _1599_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4577_ _1555_ _1566_ _1567_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3528_ _0517_ _0530_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3459_ mod.registers.r7\[8\] _2168_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3855__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _0019_ net50 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3607__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2825__I _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5274__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4583__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3394__I0 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3605__B _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4099__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ _2127_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout145_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4023__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__B _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2761_ _1638_ _2081_ _2084_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4500_ _1423_ _1462_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2692_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_8_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4326__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4362_ _0944_ _0964_ _1322_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2888__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3313_ mod.pc_2\[5\] _2432_ _0319_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4293_ _1302_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3244_ _2273_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5147__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3175_ _2191_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3065__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4262__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5297__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__I _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4014__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2959_ _2239_ _2188_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4629_ _1547_ _1371_ _1576_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3828__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__I0 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3386__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2567__A1 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4945__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_230 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3295__A2 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4492__A1 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_241 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_252 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4492__B2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_263 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_274 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_285 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_296 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4881__S _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4244__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3047__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _1793_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ _0934_ _0940_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _0857_ _0868_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4547__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2813_ _2113_ _0000_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3793_ _0683_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2744_ _2074_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ _1437_ _1823_ _2010_ mod.instr\[17\] _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4414_ _1364_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _1296_ _0590_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4276_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3227_ _2512_ _2514_ _2522_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_39_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3286__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3158_ _2427_ _2430_ _2438_ _2433_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3089_ mod.registers.r1\[0\] _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A2 _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4538__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5312__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4710__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3277__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5018__A3 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3029__A2 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4226__A1 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3201__A2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4876__S _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4130_ _0970_ _1140_ _2354_ _0512_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4061_ _1071_ _1048_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4465__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3012_ _2309_ _2278_ _2283_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _1447_ _1839_ _1835_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3914_ _0637_ _0918_ _0922_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4894_ _1657_ _1774_ _1792_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3845_ _0719_ _0824_ _0847_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3776_ _0550_ _0784_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2727_ _2063_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2951__A1 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ _2154_ _2023_ _2019_ mod.instr\[10\] _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2589_ _1853_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout102 net133 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4328_ _1289_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xfanout135 net137 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout146 net149 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4259_ _2444_ _1268_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3259__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4456__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2833__I mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3431__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3982__A3 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4144__B1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3498__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4447__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5208__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5358__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3422__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3630_ _2125_ _0639_ _0640_ _2187_ _2375_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__3574__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3561_ _0497_ _0570_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _0187_ net104 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2784__I1 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3492_ _0477_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5231_ _0118_ net99 mod.pc_1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ _0052_ net69 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4113_ _0658_ _0684_ _0851_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2918__I _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5093_ mod.instr\[4\] _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _0807_ _0984_ _0985_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_37_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout40_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2653__I _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4946_ _1456_ _1828_ _1829_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4610__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3413__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2621__B1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4877_ _1783_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3828_ _2386_ _2389_ _2399_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3759_ _0761_ _0769_ _0706_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2828__I _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4429__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3101__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2764__S _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2563__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__A3 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3340__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5114__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4953__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _1718_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2992_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4731_ _2381_ _1690_ _1692_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2603__B1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _1328_ _1585_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3159__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3613_ _0620_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3518__B _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4593_ _1523_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3544_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3475_ _2356_ _0480_ _0485_ _2342_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__4659__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4203__S0 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5214_ _0000_ _0004_ net146 mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_69_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4123__A3 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout88_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5145_ _0035_ net67 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__C _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _1930_ _1934_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ _1030_ _1037_ _0961_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4831__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2693__I0 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4929_ mod.pc_1\[0\] _1808_ _1802_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3945__I0 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3570__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2558__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5075__A1 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3389__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__I _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4889__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3561__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A3 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3260_ _0269_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3313__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3313__B2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3191_ _2488_ _2289_ _2295_ mod.registers.r4\[2\] _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5066__A1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2975_ _2256_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4041__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2931__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4714_ _1624_ _1679_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4645_ _1545_ _1426_ _1575_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ mod.registers.r1\[3\] _1561_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3527_ _2308_ _2354_ _0512_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3458_ mod.registers.r6\[8\] _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3304__A1 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__S _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3389_ _2474_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0018_ net47 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__A1 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4593__I _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5059_ _1915_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4804__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3002__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3138__A4 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3394__I1 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4099__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5048__A1 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4271__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2760_ mod.registers.r7\[12\] _2082_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout138_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2585__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2691_ mod.des.des_counter\[2\] mod.des.des_counter\[1\] mod.des.des_counter\[0\]
+ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _2238_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3129__A4 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3534__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _1359_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3582__I _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3312_ _2299_ _0320_ _0321_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ _0652_ _1197_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3243_ _2377_ _2534_ _2540_ _2341_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__A2 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ _2465_ _2467_ _2406_ _2468_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_27_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__B _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4346__C _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4262__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4014__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2958_ _2255_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2576__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2889_ _2131_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2981__C1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4628_ _1373_ _1544_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4559_ _1524_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3828__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__I1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2836__I _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5241__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3667__I _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4005__A2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_220 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_231 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_242 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3295__A3 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_253 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_264 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_275 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_286 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_297 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4244__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3930_ _0933_ _0934_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ _0584_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2812_ mod.des.des_counter\[0\] _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3792_ _0597_ _0635_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2743_ _1580_ mod.registers.r7\[5\] _2066_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2802__I0 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2674_ _2032_ _2035_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3507__A1 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4413_ mod.pc\[4\] _1365_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4344_ _1343_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _1251_ _1282_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5264__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout70_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3226_ _2523_ _2258_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3157_ _2445_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3088_ _2381_ _2382_ _2384_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4794__I0 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4171__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__I _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4474__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2566__I mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3029__A3 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5137__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5287__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4060_ _0582_ _0862_ _0870_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4465__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3011_ _2259_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4217__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ mod.pc_1\[12\] _1833_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3976__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3913_ _0794_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4893_ mod.registers.r6\[15\] _1784_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3844_ _0772_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3728__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3775_ _0785_ _0580_ _0549_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2726_ mod.des.des_dout\[15\] net11 _2059_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2657_ _1988_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4153__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _0263_ net144 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2588_ _1985_ _1295_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout103 net105 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3900__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__I _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ mod.pc0\[8\] _1319_ _1334_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xfanout114 net115 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout125 net131 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout136 net138 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout147 net149 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ mod.pc_2\[1\] _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3259__A3 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3209_ _2501_ _2189_ _2506_ _2187_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _1197_ _0813_ _1137_ _1192_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_43_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__A2 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__B2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4447__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3422__A3 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout120_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ _0495_ _0569_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ _0437_ _0464_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _0117_ net121 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _0051_ net69 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3590__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ _0777_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ _1945_ _1937_ _1946_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4438__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _0850_ _1053_ _0935_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3661__A3 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5302__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3949__B2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4945_ _1794_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3413__A3 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__A1 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4876_ _1601_ mod.registers.r6\[7\] _1770_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2621__B2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4749__I0 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3827_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3758_ _0768_ _0701_ _0710_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2709_ _2053_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3689_ _0490_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4126__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2688__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _0246_ net142 mod.des.des_dout\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4429__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2844__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2860__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2780__S _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__C _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3340__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5325__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4840__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2991_ _2161_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _1540_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2603__A1 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2603__B2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4661_ _1463_ _1556_ _1605_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3612_ _0621_ _0579_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3543_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4108__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3474_ _0481_ _0482_ _0483_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4659__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__B _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4203__S1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _0103_ net77 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4123__A4 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3331__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5144_ _0034_ net55 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5075_ mod.valid2 _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4026_ _0978_ _1010_ _1033_ _0636_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3095__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2693__I1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ mod.pc\[0\] _1806_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4859_ _1768_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3945__I1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3570__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2839__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3873__A3 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3086__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4889__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3010__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2749__I _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A4 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3313__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4510__A1 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3190_ _2286_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__B1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2974_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4713_ _0388_ _1674_ _1681_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _1438_ _1529_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3526_ _0534_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3457_ _0466_ _2316_ _2320_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3304__A2 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__A1 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3388_ _0397_ _0398_ _0390_ mod.registers.r4\[9\] _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5127_ _0017_ net50 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5057__A2 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3068__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _1470_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4009_ _1006_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3240__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5170__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4740__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2569__I mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2806__A1 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3782__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2690_ _2042_ _2039_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4731__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1248_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3311_ _2140_ _2315_ _2155_ mod.registers.r1\[5\] _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _1172_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3242_ _2535_ _2537_ _2538_ _2539_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_98_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__A3 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3173_ _2469_ _2470_ _2232_ mod.registers.r6\[2\] _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4798__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3065__A4 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3470__A1 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3222__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2957_ mod.instr_2\[2\] _2127_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5193__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2888_ _2137_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2981__B1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2981__C2 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ mod.des.des_dout\[27\] _1573_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4558_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3509_ mod.registers.r6\[14\] _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4489_ _1488_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3828__A3 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3948__I _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3461__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2852__I _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_210 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_221 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_232 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_243 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_254 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_265 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_276 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_287 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_298 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3452__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout150_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3860_ _0869_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2811_ mod.des.des_counter\[1\] _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3204__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3791_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4952__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2742_ _1570_ _2068_ _2073_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2802__I1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3593__I _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2673_ _2243_ _2030_ _2010_ mod.instr\[16\] _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4412_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4704__A1 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ _1348_ _1349_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _1283_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2937__I _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3225_ mod.pc_2\[3\] _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3156_ _2356_ _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3691__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3087_ mod.registers.r4\[0\] _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3768__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3989_ _0900_ _0327_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4794__I1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3717__B _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4599__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4548__B _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3682__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3434__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2582__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4934__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__I0 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4302__I _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2757__I _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3010_ _2268_ _2278_ _2283_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_49_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3673__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2720__I0 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4972__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2693__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3425__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4961_ _1837_ _1838_ _1835_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3912_ _0626_ _0919_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4892_ _0520_ _1773_ _1791_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ _0534_ _0850_ _0853_ _0535_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3728__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3774_ _0601_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2787__I0 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2725_ _2062_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5231__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2656_ _2017_ _2024_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4153__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2587_ _1986_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5375_ _0262_ net145 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout104 net105 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4326_ _1291_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout115 net116 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout126 net127 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout137 net138 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout148 net149 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4257_ _0531_ _2453_ _0296_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3208_ _2502_ _2503_ _2504_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4188_ _1195_ _1193_ _1198_ _0738_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2711__I0 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3139_ _2167_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2778__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4144__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2778__S _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3655__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2702__I0 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3422__A4 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5254__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4383__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3490_ _0496_ _0498_ _0500_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4967__I mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _0050_ net57 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3894__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ _0630_ _1117_ _0918_ _0977_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5091_ mod.des.des_dout\[3\] _1940_ _1941_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _0708_ _0802_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__A2 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4944_ mod.pc_1\[5\] _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4071__A1 _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3413__A4 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4875_ _1782_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2621__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3826_ _0779_ _0826_ _2448_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4749__I1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ _0689_ _0697_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2708_ mod.des.des_dout\[7\] net3 _2049_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3688_ _0698_ _0465_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4126__A2 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _1227_ _1808_ _2011_ mod.instr\[3\] _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3714__C _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5358_ _0245_ net76 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2688__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5289_ _0176_ net118 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5127__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3730__B _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2860__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5277__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4787__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3340__A3 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3628__A1 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2990_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3866__I _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2603__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3800__B2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2770__I _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4660_ _1536_ _1462_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3611_ _2525_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _1574_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3542_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4108__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3473_ _0440_ _0398_ _2418_ mod.registers.r1\[8\] _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ _0102_ net71 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _0033_ net56 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4025_ _1034_ _1035_ _0921_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2945__I mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3095__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4292__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4927_ _2190_ _1799_ _1816_ _1815_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4858_ _1771_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3809_ _0648_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4789_ _1729_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3016__I mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2855__I _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3086__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4283__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2791__S _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2597__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3010__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4310__I _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3849__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4510__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4274__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4980__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4026__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4026__B2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3596__I mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2973_ _2124_ mod.instr_2\[0\] mod.instr_2\[1\] _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4712_ _1616_ _1679_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4329__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _1519_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ mod.des.des_dout\[21\] _1543_ _1563_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3525_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2760__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ mod.registers.r5\[8\] _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3304__A3 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3387_ _2212_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5126_ _0016_ net54 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ mod.pc\[13\] _1347_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3068__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _1013_ _1017_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4017__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3240__A2 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4740__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__B _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4256__A1 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4008__A1 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3231__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2742__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3310_ _2383_ _2315_ _2291_ mod.registers.r5\[5\] _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4290_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3241_ _2211_ _2205_ _2475_ mod.registers.r1\[7\] _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3172_ _2194_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4247__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4215__I _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2956_ mod.funct3\[1\] _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3222__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2887_ _2159_ _2165_ _2170_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__2981__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _0466_ _1525_ _1611_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2981__B2 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ mod.des.des_dout\[19\] _1543_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_116_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3508_ mod.registers.r3\[14\] _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4488_ _1412_ _1489_ _1360_ _2120_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3439_ _2455_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _1936_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3461__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_200 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_211 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_222 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_233 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_244 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4229__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_255 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_266 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_277 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_288 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_299 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3452__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2810_ _2112_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout143_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3790_ _0648_ _2261_ _0649_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3204__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2741_ mod.registers.r7\[4\] _2069_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ _2032_ _2034_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4411_ _1283_ _1415_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4342_ mod.pc\[1\] _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4273_ _0774_ _1191_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4468__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3224_ _2516_ _2518_ _2520_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

