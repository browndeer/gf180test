// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire net224;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net225;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net226;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net282;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net283;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net284;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net285;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net286;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire \mod.clk ;
 wire \mod.des.des_counter[0] ;
 wire \mod.des.des_counter[1] ;
 wire \mod.des.des_counter[2] ;
 wire \mod.des.des_dout[0] ;
 wire \mod.des.des_dout[10] ;
 wire \mod.des.des_dout[11] ;
 wire \mod.des.des_dout[12] ;
 wire \mod.des.des_dout[13] ;
 wire \mod.des.des_dout[14] ;
 wire \mod.des.des_dout[15] ;
 wire \mod.des.des_dout[16] ;
 wire \mod.des.des_dout[17] ;
 wire \mod.des.des_dout[18] ;
 wire \mod.des.des_dout[19] ;
 wire \mod.des.des_dout[1] ;
 wire \mod.des.des_dout[20] ;
 wire \mod.des.des_dout[21] ;
 wire \mod.des.des_dout[22] ;
 wire \mod.des.des_dout[23] ;
 wire \mod.des.des_dout[24] ;
 wire \mod.des.des_dout[25] ;
 wire \mod.des.des_dout[26] ;
 wire \mod.des.des_dout[27] ;
 wire \mod.des.des_dout[28] ;
 wire \mod.des.des_dout[29] ;
 wire \mod.des.des_dout[2] ;
 wire \mod.des.des_dout[30] ;
 wire \mod.des.des_dout[31] ;
 wire \mod.des.des_dout[32] ;
 wire \mod.des.des_dout[33] ;
 wire \mod.des.des_dout[34] ;
 wire \mod.des.des_dout[35] ;
 wire \mod.des.des_dout[36] ;
 wire \mod.des.des_dout[3] ;
 wire \mod.des.des_dout[4] ;
 wire \mod.des.des_dout[5] ;
 wire \mod.des.des_dout[6] ;
 wire \mod.des.des_dout[7] ;
 wire \mod.des.des_dout[8] ;
 wire \mod.des.des_dout[9] ;
 wire \mod.funct3[0] ;
 wire \mod.funct3[1] ;
 wire \mod.funct3[2] ;
 wire \mod.funct7[0] ;
 wire \mod.funct7[1] ;
 wire \mod.funct7[2] ;
 wire \mod.ins_ldr_3 ;
 wire \mod.instr[0] ;
 wire \mod.instr[10] ;
 wire \mod.instr[11] ;
 wire \mod.instr[12] ;
 wire \mod.instr[13] ;
 wire \mod.instr[14] ;
 wire \mod.instr[15] ;
 wire \mod.instr[16] ;
 wire \mod.instr[17] ;
 wire \mod.instr[18] ;
 wire \mod.instr[19] ;
 wire \mod.instr[1] ;
 wire \mod.instr[20] ;
 wire \mod.instr[2] ;
 wire \mod.instr[3] ;
 wire \mod.instr[4] ;
 wire \mod.instr[5] ;
 wire \mod.instr[6] ;
 wire \mod.instr[7] ;
 wire \mod.instr[8] ;
 wire \mod.instr[9] ;
 wire \mod.instr_2[0] ;
 wire \mod.instr_2[10] ;
 wire \mod.instr_2[11] ;
 wire \mod.instr_2[12] ;
 wire \mod.instr_2[13] ;
 wire \mod.instr_2[14] ;
 wire \mod.instr_2[15] ;
 wire \mod.instr_2[16] ;
 wire \mod.instr_2[17] ;
 wire \mod.instr_2[1] ;
 wire \mod.instr_2[2] ;
 wire \mod.instr_2[3] ;
 wire \mod.instr_2[4] ;
 wire \mod.instr_2[5] ;
 wire \mod.instr_2[6] ;
 wire \mod.ldr_hzd[0] ;
 wire \mod.ldr_hzd[10] ;
 wire \mod.ldr_hzd[11] ;
 wire \mod.ldr_hzd[12] ;
 wire \mod.ldr_hzd[13] ;
 wire \mod.ldr_hzd[14] ;
 wire \mod.ldr_hzd[15] ;
 wire \mod.ldr_hzd[1] ;
 wire \mod.ldr_hzd[2] ;
 wire \mod.ldr_hzd[3] ;
 wire \mod.ldr_hzd[4] ;
 wire \mod.ldr_hzd[5] ;
 wire \mod.ldr_hzd[6] ;
 wire \mod.ldr_hzd[7] ;
 wire \mod.ldr_hzd[8] ;
 wire \mod.ldr_hzd[9] ;
 wire \mod.pc0[0] ;
 wire \mod.pc0[10] ;
 wire \mod.pc0[11] ;
 wire \mod.pc0[12] ;
 wire \mod.pc0[13] ;
 wire \mod.pc0[1] ;
 wire \mod.pc0[2] ;
 wire \mod.pc0[3] ;
 wire \mod.pc0[4] ;
 wire \mod.pc0[5] ;
 wire \mod.pc0[6] ;
 wire \mod.pc0[7] ;
 wire \mod.pc0[8] ;
 wire \mod.pc0[9] ;
 wire \mod.pc[0] ;
 wire \mod.pc[10] ;
 wire \mod.pc[11] ;
 wire \mod.pc[12] ;
 wire \mod.pc[13] ;
 wire \mod.pc[1] ;
 wire \mod.pc[2] ;
 wire \mod.pc[3] ;
 wire \mod.pc[4] ;
 wire \mod.pc[5] ;
 wire \mod.pc[6] ;
 wire \mod.pc[7] ;
 wire \mod.pc[8] ;
 wire \mod.pc[9] ;
 wire \mod.pc_1[0] ;
 wire \mod.pc_1[10] ;
 wire \mod.pc_1[11] ;
 wire \mod.pc_1[12] ;
 wire \mod.pc_1[13] ;
 wire \mod.pc_1[1] ;
 wire \mod.pc_1[2] ;
 wire \mod.pc_1[3] ;
 wire \mod.pc_1[4] ;
 wire \mod.pc_1[5] ;
 wire \mod.pc_1[6] ;
 wire \mod.pc_1[7] ;
 wire \mod.pc_1[8] ;
 wire \mod.pc_1[9] ;
 wire \mod.pc_2[0] ;
 wire \mod.pc_2[10] ;
 wire \mod.pc_2[11] ;
 wire \mod.pc_2[12] ;
 wire \mod.pc_2[13] ;
 wire \mod.pc_2[1] ;
 wire \mod.pc_2[2] ;
 wire \mod.pc_2[3] ;
 wire \mod.pc_2[4] ;
 wire \mod.pc_2[5] ;
 wire \mod.pc_2[6] ;
 wire \mod.pc_2[7] ;
 wire \mod.pc_2[8] ;
 wire \mod.pc_2[9] ;
 wire \mod.rd_3[0] ;
 wire \mod.rd_3[1] ;
 wire \mod.rd_3[2] ;
 wire \mod.rd_3[3] ;
 wire \mod.registers.r10[0] ;
 wire \mod.registers.r10[10] ;
 wire \mod.registers.r10[11] ;
 wire \mod.registers.r10[12] ;
 wire \mod.registers.r10[13] ;
 wire \mod.registers.r10[14] ;
 wire \mod.registers.r10[15] ;
 wire \mod.registers.r10[1] ;
 wire \mod.registers.r10[2] ;
 wire \mod.registers.r10[3] ;
 wire \mod.registers.r10[4] ;
 wire \mod.registers.r10[5] ;
 wire \mod.registers.r10[6] ;
 wire \mod.registers.r10[7] ;
 wire \mod.registers.r10[8] ;
 wire \mod.registers.r10[9] ;
 wire \mod.registers.r11[0] ;
 wire \mod.registers.r11[10] ;
 wire \mod.registers.r11[11] ;
 wire \mod.registers.r11[12] ;
 wire \mod.registers.r11[13] ;
 wire \mod.registers.r11[14] ;
 wire \mod.registers.r11[15] ;
 wire \mod.registers.r11[1] ;
 wire \mod.registers.r11[2] ;
 wire \mod.registers.r11[3] ;
 wire \mod.registers.r11[4] ;
 wire \mod.registers.r11[5] ;
 wire \mod.registers.r11[6] ;
 wire \mod.registers.r11[7] ;
 wire \mod.registers.r11[8] ;
 wire \mod.registers.r11[9] ;
 wire \mod.registers.r12[0] ;
 wire \mod.registers.r12[10] ;
 wire \mod.registers.r12[11] ;
 wire \mod.registers.r12[12] ;
 wire \mod.registers.r12[13] ;
 wire \mod.registers.r12[14] ;
 wire \mod.registers.r12[15] ;
 wire \mod.registers.r12[1] ;
 wire \mod.registers.r12[2] ;
 wire \mod.registers.r12[3] ;
 wire \mod.registers.r12[4] ;
 wire \mod.registers.r12[5] ;
 wire \mod.registers.r12[6] ;
 wire \mod.registers.r12[7] ;
 wire \mod.registers.r12[8] ;
 wire \mod.registers.r12[9] ;
 wire \mod.registers.r13[0] ;
 wire \mod.registers.r13[10] ;
 wire \mod.registers.r13[11] ;
 wire \mod.registers.r13[12] ;
 wire \mod.registers.r13[13] ;
 wire \mod.registers.r13[14] ;
 wire \mod.registers.r13[15] ;
 wire \mod.registers.r13[1] ;
 wire \mod.registers.r13[2] ;
 wire \mod.registers.r13[3] ;
 wire \mod.registers.r13[4] ;
 wire \mod.registers.r13[5] ;
 wire \mod.registers.r13[6] ;
 wire \mod.registers.r13[7] ;
 wire \mod.registers.r13[8] ;
 wire \mod.registers.r13[9] ;
 wire \mod.registers.r14[0] ;
 wire \mod.registers.r14[10] ;
 wire \mod.registers.r14[11] ;
 wire \mod.registers.r14[12] ;
 wire \mod.registers.r14[13] ;
 wire \mod.registers.r14[14] ;
 wire \mod.registers.r14[15] ;
 wire \mod.registers.r14[1] ;
 wire \mod.registers.r14[2] ;
 wire \mod.registers.r14[3] ;
 wire \mod.registers.r14[4] ;
 wire \mod.registers.r14[5] ;
 wire \mod.registers.r14[6] ;
 wire \mod.registers.r14[7] ;
 wire \mod.registers.r14[8] ;
 wire \mod.registers.r14[9] ;
 wire \mod.registers.r15[0] ;
 wire \mod.registers.r15[10] ;
 wire \mod.registers.r15[11] ;
 wire \mod.registers.r15[12] ;
 wire \mod.registers.r15[13] ;
 wire \mod.registers.r15[14] ;
 wire \mod.registers.r15[15] ;
 wire \mod.registers.r15[1] ;
 wire \mod.registers.r15[2] ;
 wire \mod.registers.r15[3] ;
 wire \mod.registers.r15[4] ;
 wire \mod.registers.r15[5] ;
 wire \mod.registers.r15[6] ;
 wire \mod.registers.r15[7] ;
 wire \mod.registers.r15[8] ;
 wire \mod.registers.r15[9] ;
 wire \mod.registers.r1[0] ;
 wire \mod.registers.r1[10] ;
 wire \mod.registers.r1[11] ;
 wire \mod.registers.r1[12] ;
 wire \mod.registers.r1[13] ;
 wire \mod.registers.r1[14] ;
 wire \mod.registers.r1[15] ;
 wire \mod.registers.r1[1] ;
 wire \mod.registers.r1[2] ;
 wire \mod.registers.r1[3] ;
 wire \mod.registers.r1[4] ;
 wire \mod.registers.r1[5] ;
 wire \mod.registers.r1[6] ;
 wire \mod.registers.r1[7] ;
 wire \mod.registers.r1[8] ;
 wire \mod.registers.r1[9] ;
 wire \mod.registers.r2[0] ;
 wire \mod.registers.r2[10] ;
 wire \mod.registers.r2[11] ;
 wire \mod.registers.r2[12] ;
 wire \mod.registers.r2[13] ;
 wire \mod.registers.r2[14] ;
 wire \mod.registers.r2[15] ;
 wire \mod.registers.r2[1] ;
 wire \mod.registers.r2[2] ;
 wire \mod.registers.r2[3] ;
 wire \mod.registers.r2[4] ;
 wire \mod.registers.r2[5] ;
 wire \mod.registers.r2[6] ;
 wire \mod.registers.r2[7] ;
 wire \mod.registers.r2[8] ;
 wire \mod.registers.r2[9] ;
 wire \mod.registers.r3[0] ;
 wire \mod.registers.r3[10] ;
 wire \mod.registers.r3[11] ;
 wire \mod.registers.r3[12] ;
 wire \mod.registers.r3[13] ;
 wire \mod.registers.r3[14] ;
 wire \mod.registers.r3[15] ;
 wire \mod.registers.r3[1] ;
 wire \mod.registers.r3[2] ;
 wire \mod.registers.r3[3] ;
 wire \mod.registers.r3[4] ;
 wire \mod.registers.r3[5] ;
 wire \mod.registers.r3[6] ;
 wire \mod.registers.r3[7] ;
 wire \mod.registers.r3[8] ;
 wire \mod.registers.r3[9] ;
 wire \mod.registers.r4[0] ;
 wire \mod.registers.r4[10] ;
 wire \mod.registers.r4[11] ;
 wire \mod.registers.r4[12] ;
 wire \mod.registers.r4[13] ;
 wire \mod.registers.r4[14] ;
 wire \mod.registers.r4[15] ;
 wire \mod.registers.r4[1] ;
 wire \mod.registers.r4[2] ;
 wire \mod.registers.r4[3] ;
 wire \mod.registers.r4[4] ;
 wire \mod.registers.r4[5] ;
 wire \mod.registers.r4[6] ;
 wire \mod.registers.r4[7] ;
 wire \mod.registers.r4[8] ;
 wire \mod.registers.r4[9] ;
 wire \mod.registers.r5[0] ;
 wire \mod.registers.r5[10] ;
 wire \mod.registers.r5[11] ;
 wire \mod.registers.r5[12] ;
 wire \mod.registers.r5[13] ;
 wire \mod.registers.r5[14] ;
 wire \mod.registers.r5[15] ;
 wire \mod.registers.r5[1] ;
 wire \mod.registers.r5[2] ;
 wire \mod.registers.r5[3] ;
 wire \mod.registers.r5[4] ;
 wire \mod.registers.r5[5] ;
 wire \mod.registers.r5[6] ;
 wire \mod.registers.r5[7] ;
 wire \mod.registers.r5[8] ;
 wire \mod.registers.r5[9] ;
 wire \mod.registers.r6[0] ;
 wire \mod.registers.r6[10] ;
 wire \mod.registers.r6[11] ;
 wire \mod.registers.r6[12] ;
 wire \mod.registers.r6[13] ;
 wire \mod.registers.r6[14] ;
 wire \mod.registers.r6[15] ;
 wire \mod.registers.r6[1] ;
 wire \mod.registers.r6[2] ;
 wire \mod.registers.r6[3] ;
 wire \mod.registers.r6[4] ;
 wire \mod.registers.r6[5] ;
 wire \mod.registers.r6[6] ;
 wire \mod.registers.r6[7] ;
 wire \mod.registers.r6[8] ;
 wire \mod.registers.r6[9] ;
 wire \mod.registers.r7[0] ;
 wire \mod.registers.r7[10] ;
 wire \mod.registers.r7[11] ;
 wire \mod.registers.r7[12] ;
 wire \mod.registers.r7[13] ;
 wire \mod.registers.r7[14] ;
 wire \mod.registers.r7[15] ;
 wire \mod.registers.r7[1] ;
 wire \mod.registers.r7[2] ;
 wire \mod.registers.r7[3] ;
 wire \mod.registers.r7[4] ;
 wire \mod.registers.r7[5] ;
 wire \mod.registers.r7[6] ;
 wire \mod.registers.r7[7] ;
 wire \mod.registers.r7[8] ;
 wire \mod.registers.r7[9] ;
 wire \mod.registers.r8[0] ;
 wire \mod.registers.r8[10] ;
 wire \mod.registers.r8[11] ;
 wire \mod.registers.r8[12] ;
 wire \mod.registers.r8[13] ;
 wire \mod.registers.r8[14] ;
 wire \mod.registers.r8[15] ;
 wire \mod.registers.r8[1] ;
 wire \mod.registers.r8[2] ;
 wire \mod.registers.r8[3] ;
 wire \mod.registers.r8[4] ;
 wire \mod.registers.r8[5] ;
 wire \mod.registers.r8[6] ;
 wire \mod.registers.r8[7] ;
 wire \mod.registers.r8[8] ;
 wire \mod.registers.r8[9] ;
 wire \mod.registers.r9[0] ;
 wire \mod.registers.r9[10] ;
 wire \mod.registers.r9[11] ;
 wire \mod.registers.r9[12] ;
 wire \mod.registers.r9[13] ;
 wire \mod.registers.r9[14] ;
 wire \mod.registers.r9[15] ;
 wire \mod.registers.r9[1] ;
 wire \mod.registers.r9[2] ;
 wire \mod.registers.r9[3] ;
 wire \mod.registers.r9[4] ;
 wire \mod.registers.r9[5] ;
 wire \mod.registers.r9[6] ;
 wire \mod.registers.r9[7] ;
 wire \mod.registers.r9[8] ;
 wire \mod.registers.r9[9] ;
 wire \mod.ri_3 ;
 wire \mod.valid0 ;
 wire \mod.valid1 ;
 wire \mod.valid2 ;
 wire \mod.valid_out3 ;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net350;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net351;
 wire net379;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3293_ (.I(\mod.des.des_counter[0] ),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3294_ (.I(\mod.des.des_counter[1] ),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3295_ (.A1(_0000_),
    .A2(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3296_ (.A1(net176),
    .A2(_3151_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3297_ (.I(_3152_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3298_ (.A1(\mod.des.des_counter[0] ),
    .A2(_3150_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3299_ (.A1(_0000_),
    .A2(\mod.des.des_counter[1] ),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3300_ (.A1(_3153_),
    .A2(_3154_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3301_ (.I(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3302_ (.I(_3156_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3303_ (.A1(\mod.des.des_counter[2] ),
    .A2(_3151_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3304_ (.I(_3157_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3305_ (.I(\mod.instr_2[15] ),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3306_ (.I(\mod.instr_2[14] ),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3307_ (.A1(_3158_),
    .A2(_3159_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3308_ (.I(\mod.instr_2[17] ),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3309_ (.I(\mod.instr_2[16] ),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3310_ (.A1(_3161_),
    .A2(_3162_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3311_ (.A1(_3160_),
    .A2(_3163_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3312_ (.I(_3164_),
    .Z(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3313_ (.I(_3161_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3314_ (.I(\mod.instr_2[16] ),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3315_ (.I(_3167_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3316_ (.A1(_3166_),
    .A2(_3168_),
    .A3(_3160_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3317_ (.I(_3169_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3318_ (.A1(\mod.registers.r3[0] ),
    .A2(_3165_),
    .B1(_3170_),
    .B2(\mod.registers.r7[0] ),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3319_ (.A1(_3158_),
    .A2(_3159_),
    .Z(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3320_ (.A1(_3166_),
    .A2(_3168_),
    .A3(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3321_ (.I(_3173_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3322_ (.I(\mod.instr_2[15] ),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3323_ (.I(\mod.instr_2[14] ),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3324_ (.A1(_3175_),
    .A2(_3176_),
    .A3(_3163_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3325_ (.I(_3177_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3326_ (.A1(\mod.registers.r4[0] ),
    .A2(_3174_),
    .B1(_3178_),
    .B2(\mod.registers.r1[0] ),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3327_ (.A1(_3171_),
    .A2(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3328_ (.I(_3161_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3329_ (.I(\mod.instr_2[15] ),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3330_ (.I(_3182_),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3331_ (.I(\mod.instr_2[14] ),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3332_ (.A1(_3181_),
    .A2(_3167_),
    .A3(_3183_),
    .A4(_3184_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3333_ (.I(_3185_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3334_ (.I(_3176_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3335_ (.A1(_3166_),
    .A2(_3167_),
    .A3(_3175_),
    .A4(_3187_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3336_ (.I(_3188_),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3337_ (.A1(_3182_),
    .A2(_3159_),
    .A3(_3163_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3338_ (.I(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3339_ (.A1(\mod.registers.r6[0] ),
    .A2(_3186_),
    .B1(_3189_),
    .B2(\mod.registers.r5[0] ),
    .C1(\mod.registers.r2[0] ),
    .C2(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3340_ (.I(\mod.instr_2[17] ),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3341_ (.A1(_3193_),
    .A2(_3162_),
    .A3(_3182_),
    .A4(_3184_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3342_ (.I(_3194_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3343_ (.I(_3193_),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3344_ (.I(\mod.instr_2[16] ),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3345_ (.A1(_3196_),
    .A2(_3197_),
    .A3(_3175_),
    .A4(_3187_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3346_ (.I(_3198_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3347_ (.A1(\mod.registers.r10[0] ),
    .A2(_3195_),
    .B1(_3199_),
    .B2(\mod.registers.r9[0] ),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3348_ (.A1(_3196_),
    .A2(_3197_),
    .A3(_3160_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3349_ (.I(_3201_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3350_ (.A1(_3196_),
    .A2(_3197_),
    .A3(_3172_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3351_ (.I(_3203_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3352_ (.A1(\mod.registers.r11[0] ),
    .A2(_3202_),
    .B1(_3204_),
    .B2(\mod.registers.r8[0] ),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3353_ (.A1(_3161_),
    .A2(\mod.instr_2[16] ),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3354_ (.A1(_3183_),
    .A2(_3184_),
    .A3(_3206_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3355_ (.I(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3356_ (.I(_3158_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3357_ (.A1(_3209_),
    .A2(_3187_),
    .A3(_3206_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3358_ (.I(_3210_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3359_ (.I(\mod.registers.r12[0] ),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3360_ (.I(_3172_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3361_ (.I(_3206_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3362_ (.I(_3181_),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3363_ (.I(_3162_),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3364_ (.I(_3159_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3365_ (.A1(_3215_),
    .A2(_3216_),
    .A3(_3209_),
    .A4(_3217_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3366_ (.I(\mod.registers.r15[0] ),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3367_ (.A1(_3212_),
    .A2(_3213_),
    .A3(_3214_),
    .B1(_3218_),
    .B2(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3368_ (.A1(\mod.registers.r14[0] ),
    .A2(_3208_),
    .B1(_3211_),
    .B2(\mod.registers.r13[0] ),
    .C(_3220_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3369_ (.A1(_3192_),
    .A2(_3200_),
    .A3(_3205_),
    .A4(_3221_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3370_ (.I(_3153_),
    .Z(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3371_ (.A1(_3180_),
    .A2(_3222_),
    .B(_3223_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3372_ (.I(_3154_),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3373_ (.I(\mod.funct3[2] ),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3374_ (.I(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3375_ (.I(\mod.funct3[1] ),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3376_ (.I(_3228_),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3377_ (.I(\mod.instr_2[2] ),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3378_ (.I(\mod.instr_2[0] ),
    .Z(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3379_ (.A1(_3230_),
    .A2(_3231_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3380_ (.I(_3232_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3381_ (.I(\mod.instr_2[1] ),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3382_ (.A1(_3230_),
    .A2(_3231_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3383_ (.A1(_3234_),
    .A2(_3235_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3384_ (.I(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3385_ (.I(_3237_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3386_ (.I(_3238_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3387_ (.A1(_3233_),
    .A2(_3239_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3388_ (.A1(_3227_),
    .A2(_3229_),
    .A3(_3240_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3389_ (.I(_3241_),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3390_ (.I(_3242_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3391_ (.I(_3233_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3392_ (.I(_3238_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3393_ (.I(_3245_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3394_ (.I(_3246_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3395_ (.I(_3226_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3396_ (.A1(_3248_),
    .A2(_3228_),
    .A3(\mod.funct3[0] ),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3397_ (.A1(_3244_),
    .A2(_3247_),
    .A3(_3249_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3398_ (.A1(_3230_),
    .A2(_3231_),
    .B(\mod.instr_2[1] ),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3399_ (.I(_3251_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3400_ (.I(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3401_ (.I(_3252_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3402_ (.I(\mod.instr_2[3] ),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3403_ (.I(_3187_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3404_ (.A1(\mod.instr_2[2] ),
    .A2(\mod.instr_2[0] ),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3405_ (.A1(\mod.funct3[2] ),
    .A2(_3232_),
    .B(_3257_),
    .C(_3234_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3406_ (.I0(_3255_),
    .I1(_3256_),
    .S(_3258_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3407_ (.A1(_3254_),
    .A2(_3259_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3408_ (.A1(_3253_),
    .A2(_3180_),
    .A3(_3222_),
    .B(_3260_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3409_ (.I(_3261_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3410_ (.I(\mod.pc_2[0] ),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3411_ (.I(_3236_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3412_ (.I(_3264_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3413_ (.I(_3265_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3414_ (.I(\mod.instr_2[13] ),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3415_ (.I(\mod.instr_2[12] ),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3416_ (.I(_3268_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3417_ (.A1(\mod.instr_2[11] ),
    .A2(\mod.instr_2[10] ),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3418_ (.A1(_3267_),
    .A2(_3269_),
    .A3(_3270_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3419_ (.I(_3271_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3420_ (.I(_3272_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3421_ (.I(\mod.instr_2[11] ),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3422_ (.I(_3274_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3423_ (.I(\mod.instr_2[10] ),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3424_ (.I(_3276_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3425_ (.A1(_3267_),
    .A2(_3269_),
    .A3(_3275_),
    .A4(_3277_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_3278_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3427_ (.A1(\mod.registers.r8[0] ),
    .A2(_3273_),
    .B1(_3279_),
    .B2(\mod.registers.r10[0] ),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3428_ (.A1(\mod.instr_2[13] ),
    .A2(_3268_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3429_ (.A1(_3275_),
    .A2(_3277_),
    .A3(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3430_ (.I(_3282_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3431_ (.I(\mod.instr_2[13] ),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3432_ (.I(\mod.instr_2[12] ),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3433_ (.A1(_3284_),
    .A2(_3285_),
    .A3(_3274_),
    .A4(_3276_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3434_ (.I(_3286_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3435_ (.A1(\mod.registers.r14[0] ),
    .A2(_3283_),
    .B1(_3287_),
    .B2(\mod.registers.r6[0] ),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3436_ (.A1(\mod.instr_2[11] ),
    .A2(_3276_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3437_ (.A1(_3267_),
    .A2(_3269_),
    .A3(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3438_ (.I(_3290_),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3439_ (.I(_3291_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3440_ (.A1(_3284_),
    .A2(_3268_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3441_ (.A1(_3275_),
    .A2(_3277_),
    .A3(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3442_ (.I(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3443_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3444_ (.A1(\mod.registers.r11[0] ),
    .A2(_3292_),
    .B1(_0413_),
    .B2(\mod.registers.r2[0] ),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3445_ (.I(_3284_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3446_ (.I(_3285_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3447_ (.I(_3270_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3448_ (.A1(_0415_),
    .A2(_0416_),
    .A3(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3449_ (.I(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3450_ (.I(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3451_ (.I(_3236_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3452_ (.A1(\mod.registers.r4[0] ),
    .A2(_0420_),
    .B(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3453_ (.A1(_3280_),
    .A2(_3288_),
    .A3(_0414_),
    .A4(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3454_ (.I(_3267_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3455_ (.I(\mod.instr_2[11] ),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3456_ (.I(\mod.instr_2[10] ),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3457_ (.A1(_0424_),
    .A2(_3269_),
    .A3(_0425_),
    .A4(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3458_ (.I(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3459_ (.I(_3289_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3460_ (.A1(_0429_),
    .A2(_0410_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3461_ (.I(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3462_ (.A1(\mod.registers.r9[0] ),
    .A2(_0428_),
    .B1(_0431_),
    .B2(\mod.registers.r3[0] ),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3463_ (.I(_3281_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3464_ (.A1(_0429_),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3465_ (.I(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3466_ (.A1(_3281_),
    .A2(_0417_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3467_ (.I(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3468_ (.A1(\mod.registers.r15[0] ),
    .A2(_0435_),
    .B1(_0437_),
    .B2(\mod.registers.r12[0] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3469_ (.A1(_3284_),
    .A2(_0416_),
    .A3(_0425_),
    .A4(_0426_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3470_ (.I(_0439_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3471_ (.A1(_0415_),
    .A2(_0416_),
    .A3(_3289_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3472_ (.I(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3473_ (.A1(\mod.registers.r5[0] ),
    .A2(_0440_),
    .B1(_0442_),
    .B2(\mod.registers.r7[0] ),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3474_ (.I(_0425_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3475_ (.I(_0426_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3476_ (.A1(_0444_),
    .A2(_0445_),
    .A3(_3281_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3477_ (.I(_0446_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3478_ (.A1(_0444_),
    .A2(_0445_),
    .A3(_0410_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3479_ (.I(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3480_ (.A1(\mod.registers.r13[0] ),
    .A2(_0447_),
    .B1(_0449_),
    .B2(\mod.registers.r1[0] ),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3481_ (.A1(_0432_),
    .A2(_0438_),
    .A3(_0443_),
    .A4(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3482_ (.A1(_3263_),
    .A2(_3266_),
    .B1(_0423_),
    .B2(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3483_ (.I(_0452_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3484_ (.A1(_3246_),
    .A2(_3262_),
    .A3(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3485_ (.A1(_3254_),
    .A2(_3180_),
    .A3(_3222_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3486_ (.I(_3234_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3487_ (.I(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3488_ (.I(_3237_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3489_ (.A1(_0457_),
    .A2(_3259_),
    .B(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3490_ (.A1(_0455_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3491_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3492_ (.A1(_0461_),
    .A2(_0453_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3493_ (.A1(_0454_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3494_ (.I(_3265_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3495_ (.I(_3173_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3496_ (.I(_3177_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3497_ (.A1(\mod.registers.r4[1] ),
    .A2(_0465_),
    .B1(_0466_),
    .B2(\mod.registers.r1[1] ),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3498_ (.I(_3188_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3499_ (.A1(\mod.registers.r2[1] ),
    .A2(_3191_),
    .B1(_0468_),
    .B2(\mod.registers.r5[1] ),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_0467_),
    .A2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3501_ (.I(_3164_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3502_ (.A1(\mod.registers.r3[1] ),
    .A2(_0471_),
    .B1(_3186_),
    .B2(\mod.registers.r6[1] ),
    .C1(\mod.registers.r7[1] ),
    .C2(_3170_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3503_ (.I(_3203_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3504_ (.A1(\mod.registers.r8[1] ),
    .A2(_0473_),
    .B1(_3199_),
    .B2(\mod.registers.r9[1] ),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3505_ (.A1(\mod.registers.r11[1] ),
    .A2(_3202_),
    .B1(_3195_),
    .B2(\mod.registers.r10[1] ),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3506_ (.A1(_3175_),
    .A2(_3217_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3507_ (.A1(_3181_),
    .A2(_3162_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3508_ (.I(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3509_ (.A1(\mod.registers.r12[1] ),
    .A2(_0476_),
    .A3(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3510_ (.I(_3209_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3511_ (.A1(_0480_),
    .A2(_3256_),
    .A3(\mod.registers.r14[1] ),
    .A4(_0477_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3512_ (.I(_3183_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3513_ (.I(_3217_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3514_ (.A1(_0482_),
    .A2(_0483_),
    .A3(\mod.registers.r13[1] ),
    .A4(_0477_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3515_ (.A1(_3181_),
    .A2(_3197_),
    .A3(_3158_),
    .A4(_3184_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3516_ (.A1(\mod.registers.r15[1] ),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3517_ (.A1(_0479_),
    .A2(_0481_),
    .A3(_0484_),
    .A4(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3518_ (.A1(_0472_),
    .A2(_0474_),
    .A3(_0475_),
    .A4(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3519_ (.I(_3252_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3520_ (.I(\mod.instr_2[4] ),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3521_ (.I0(_0490_),
    .I1(_0482_),
    .S(_3258_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3522_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3523_ (.A1(_0489_),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3524_ (.A1(_3254_),
    .A2(_0470_),
    .A3(_0488_),
    .B(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3525_ (.A1(_0464_),
    .A2(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3526_ (.I(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3527_ (.I(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3528_ (.A1(_0457_),
    .A2(_3257_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3529_ (.I(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3530_ (.I(_3278_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3531_ (.A1(\mod.registers.r8[6] ),
    .A2(_3272_),
    .B1(_0500_),
    .B2(\mod.registers.r10[6] ),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3532_ (.I(_3282_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3533_ (.I(_3286_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3534_ (.A1(\mod.registers.r14[6] ),
    .A2(_0502_),
    .B1(_0503_),
    .B2(\mod.registers.r6[6] ),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3535_ (.I(_3290_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3536_ (.I(_0411_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3537_ (.A1(\mod.registers.r11[6] ),
    .A2(_0505_),
    .B1(_0506_),
    .B2(\mod.registers.r2[6] ),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3538_ (.I(_0418_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3539_ (.A1(\mod.registers.r4[6] ),
    .A2(_0508_),
    .B(_3237_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3540_ (.A1(_0501_),
    .A2(_0504_),
    .A3(_0507_),
    .A4(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3541_ (.I(_0427_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3542_ (.I(_0430_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3543_ (.A1(\mod.registers.r9[6] ),
    .A2(_0511_),
    .B1(_0512_),
    .B2(\mod.registers.r3[6] ),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3544_ (.I(_0434_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3545_ (.I(_0436_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3546_ (.A1(\mod.registers.r15[6] ),
    .A2(_0514_),
    .B1(_0515_),
    .B2(\mod.registers.r12[6] ),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3547_ (.I(_0439_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3548_ (.I(_0441_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3549_ (.A1(\mod.registers.r5[6] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\mod.registers.r7[6] ),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3550_ (.I(_0446_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3551_ (.I(_0448_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3552_ (.A1(\mod.registers.r13[6] ),
    .A2(_0520_),
    .B1(_0521_),
    .B2(\mod.registers.r1[6] ),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3553_ (.A1(_0513_),
    .A2(_0516_),
    .A3(_0519_),
    .A4(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3554_ (.A1(\mod.pc_2[6] ),
    .A2(_0499_),
    .B1(_0510_),
    .B2(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3555_ (.I(_0524_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3556_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3557_ (.I(_0460_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3558_ (.I(_0464_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3559_ (.I(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3560_ (.I(\mod.pc_2[7] ),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3561_ (.I(_3271_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3562_ (.I(_3278_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3563_ (.A1(\mod.registers.r8[7] ),
    .A2(_0531_),
    .B1(_0532_),
    .B2(\mod.registers.r10[7] ),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3564_ (.I(_3282_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3565_ (.I(_3286_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3566_ (.A1(\mod.registers.r14[7] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\mod.registers.r6[7] ),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3567_ (.A1(\mod.registers.r11[7] ),
    .A2(_0505_),
    .B1(_0506_),
    .B2(\mod.registers.r2[7] ),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3568_ (.A1(\mod.registers.r4[7] ),
    .A2(_0508_),
    .B(_3237_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3569_ (.A1(_0533_),
    .A2(_0536_),
    .A3(_0537_),
    .A4(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3570_ (.A1(\mod.registers.r15[7] ),
    .A2(_0435_),
    .B1(_0437_),
    .B2(\mod.registers.r12[7] ),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3571_ (.I(_0446_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3572_ (.I(_0448_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3573_ (.A1(\mod.registers.r13[7] ),
    .A2(_0541_),
    .B1(_0542_),
    .B2(\mod.registers.r1[7] ),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3574_ (.I(_0427_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3575_ (.I(_0430_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3576_ (.A1(\mod.registers.r9[7] ),
    .A2(_0544_),
    .B1(_0545_),
    .B2(\mod.registers.r3[7] ),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3577_ (.I(_0439_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3578_ (.I(_0441_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3579_ (.A1(\mod.registers.r5[7] ),
    .A2(_0547_),
    .B1(_0548_),
    .B2(\mod.registers.r7[7] ),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3580_ (.A1(_0540_),
    .A2(_0543_),
    .A3(_0546_),
    .A4(_0549_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3581_ (.A1(_0530_),
    .A2(_0528_),
    .B1(_0539_),
    .B2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3582_ (.I(_3261_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3583_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3584_ (.A1(_0529_),
    .A2(_0551_),
    .A3(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3585_ (.A1(_0526_),
    .A2(_0527_),
    .B(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3586_ (.I(_0455_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3587_ (.I(_0459_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3588_ (.A1(\mod.registers.r7[4] ),
    .A2(_0442_),
    .B1(_3273_),
    .B2(\mod.registers.r8[4] ),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3589_ (.A1(\mod.registers.r14[4] ),
    .A2(_3283_),
    .B1(_3287_),
    .B2(\mod.registers.r6[4] ),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3590_ (.I(_3234_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3591_ (.I(_3235_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3592_ (.I(_3268_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3593_ (.A1(_0415_),
    .A2(_0562_),
    .A3(_0444_),
    .A4(_3277_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3594_ (.I(\mod.registers.r15[4] ),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3595_ (.A1(_0560_),
    .A2(_0561_),
    .B1(_0563_),
    .B2(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3596_ (.A1(\mod.registers.r13[4] ),
    .A2(_0447_),
    .B1(_0431_),
    .B2(\mod.registers.r3[4] ),
    .C(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3597_ (.A1(_0558_),
    .A2(_0559_),
    .A3(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3598_ (.A1(\mod.registers.r10[4] ),
    .A2(_3279_),
    .B1(_0413_),
    .B2(\mod.registers.r2[4] ),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3599_ (.A1(\mod.registers.r4[4] ),
    .A2(_0420_),
    .B1(_0449_),
    .B2(\mod.registers.r1[4] ),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3600_ (.A1(\mod.registers.r12[4] ),
    .A2(_0437_),
    .B1(_0428_),
    .B2(\mod.registers.r9[4] ),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3601_ (.A1(\mod.registers.r5[4] ),
    .A2(_0440_),
    .B1(_3292_),
    .B2(\mod.registers.r11[4] ),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3602_ (.A1(_0568_),
    .A2(_0569_),
    .A3(_0570_),
    .A4(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3603_ (.A1(\mod.pc_2[4] ),
    .A2(_0499_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3604_ (.A1(_0567_),
    .A2(_0572_),
    .B(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3605_ (.A1(_0556_),
    .A2(_0557_),
    .B(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3606_ (.I(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3607_ (.I(_3265_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3608_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3609_ (.I(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3610_ (.I(\mod.pc_2[5] ),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3611_ (.A1(\mod.registers.r8[5] ),
    .A2(_3271_),
    .B1(_3278_),
    .B2(\mod.registers.r10[5] ),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3612_ (.A1(\mod.registers.r14[5] ),
    .A2(_3282_),
    .B1(_3286_),
    .B2(\mod.registers.r6[5] ),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3613_ (.A1(\mod.registers.r11[5] ),
    .A2(_3291_),
    .B1(_0411_),
    .B2(\mod.registers.r2[5] ),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3614_ (.A1(\mod.registers.r4[5] ),
    .A2(_0418_),
    .B(_3236_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3615_ (.A1(_0581_),
    .A2(_0582_),
    .A3(_0583_),
    .A4(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3616_ (.A1(\mod.registers.r15[5] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.registers.r12[5] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3617_ (.A1(\mod.registers.r9[5] ),
    .A2(_0427_),
    .B1(_0430_),
    .B2(\mod.registers.r3[5] ),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3618_ (.A1(\mod.registers.r5[5] ),
    .A2(_0439_),
    .B1(_0441_),
    .B2(\mod.registers.r7[5] ),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3619_ (.A1(\mod.registers.r13[5] ),
    .A2(_0446_),
    .B1(_0448_),
    .B2(\mod.registers.r1[5] ),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3620_ (.A1(_0586_),
    .A2(_0587_),
    .A3(_0588_),
    .A4(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3621_ (.A1(_0580_),
    .A2(_0421_),
    .B1(_0585_),
    .B2(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3622_ (.A1(_0579_),
    .A2(_0591_),
    .A3(_3262_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3623_ (.I(_0495_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3624_ (.A1(_0576_),
    .A2(_0592_),
    .B(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3625_ (.I(_0489_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3626_ (.I(_3169_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3627_ (.A1(\mod.registers.r3[2] ),
    .A2(_3165_),
    .B1(_0596_),
    .B2(\mod.registers.r7[2] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3628_ (.A1(\mod.registers.r4[2] ),
    .A2(_3174_),
    .B1(_3178_),
    .B2(\mod.registers.r1[2] ),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3629_ (.A1(_0597_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3630_ (.I(_3185_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3631_ (.A1(\mod.registers.r6[2] ),
    .A2(_0600_),
    .B1(_3189_),
    .B2(\mod.registers.r5[2] ),
    .C1(\mod.registers.r2[2] ),
    .C2(_3191_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3632_ (.I(_3194_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3633_ (.I(_3198_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3634_ (.A1(\mod.registers.r10[2] ),
    .A2(_0602_),
    .B1(_0603_),
    .B2(\mod.registers.r9[2] ),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3635_ (.I(_3201_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3636_ (.A1(\mod.registers.r11[2] ),
    .A2(_0605_),
    .B1(_0473_),
    .B2(\mod.registers.r8[2] ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3637_ (.I(_3207_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3638_ (.I(_3210_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3639_ (.I(\mod.registers.r12[2] ),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3640_ (.I(\mod.registers.r15[2] ),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3641_ (.A1(_0609_),
    .A2(_3213_),
    .A3(_3214_),
    .B1(_3218_),
    .B2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3642_ (.A1(\mod.registers.r14[2] ),
    .A2(_0607_),
    .B1(_0608_),
    .B2(\mod.registers.r13[2] ),
    .C(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3643_ (.A1(_0601_),
    .A2(_0604_),
    .A3(_0606_),
    .A4(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3644_ (.A1(_0456_),
    .A2(_3235_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3645_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3646_ (.I(_3216_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3647_ (.I(_3258_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3648_ (.I0(\mod.instr_2[5] ),
    .I1(_0616_),
    .S(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3649_ (.A1(_0615_),
    .A2(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3650_ (.A1(_0595_),
    .A2(_0599_),
    .A3(_0613_),
    .B(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3651_ (.A1(_0578_),
    .A2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3652_ (.I(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3653_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3654_ (.A1(_0497_),
    .A2(_0555_),
    .B(_0594_),
    .C(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3655_ (.I(_0495_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3656_ (.A1(_0625_),
    .A2(_0622_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3657_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3658_ (.I(\mod.pc_2[2] ),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3659_ (.A1(\mod.registers.r8[2] ),
    .A2(_0531_),
    .B1(_0532_),
    .B2(\mod.registers.r10[2] ),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3660_ (.A1(\mod.registers.r14[2] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\mod.registers.r6[2] ),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3661_ (.I(_0415_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3662_ (.I(_0416_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3663_ (.I(_3276_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3664_ (.A1(_0444_),
    .A2(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3665_ (.A1(_0631_),
    .A2(_0632_),
    .A3(\mod.registers.r11[2] ),
    .A4(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3666_ (.I(_0562_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3667_ (.I(_0425_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3668_ (.A1(_0637_),
    .A2(_0633_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3669_ (.A1(_0424_),
    .A2(_0636_),
    .A3(\mod.registers.r4[2] ),
    .A4(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3670_ (.A1(_0631_),
    .A2(_0562_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3671_ (.A1(_0637_),
    .A2(_0445_),
    .A3(\mod.registers.r2[2] ),
    .A4(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3672_ (.A1(_0498_),
    .A2(_0635_),
    .A3(_0639_),
    .A4(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3673_ (.A1(_0629_),
    .A2(_0630_),
    .A3(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3674_ (.A1(\mod.registers.r7[2] ),
    .A2(_0548_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3675_ (.A1(\mod.registers.r5[2] ),
    .A2(_0547_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3676_ (.A1(\mod.registers.r9[2] ),
    .A2(_0544_),
    .B1(_0545_),
    .B2(\mod.registers.r3[2] ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3677_ (.A1(_0609_),
    .A2(_0433_),
    .A3(_0417_),
    .B1(_0563_),
    .B2(_0610_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3678_ (.A1(\mod.registers.r13[2] ),
    .A2(_0541_),
    .B1(_0542_),
    .B2(\mod.registers.r1[2] ),
    .C(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3679_ (.A1(_0644_),
    .A2(_0645_),
    .A3(_0646_),
    .A4(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3680_ (.A1(_0628_),
    .A2(_0577_),
    .B1(_0643_),
    .B2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3681_ (.I(\mod.pc_2[3] ),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3682_ (.A1(\mod.registers.r8[3] ),
    .A2(_0531_),
    .B1(_0532_),
    .B2(\mod.registers.r10[3] ),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3683_ (.A1(\mod.registers.r14[3] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\mod.registers.r6[3] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3684_ (.A1(\mod.registers.r11[3] ),
    .A2(_0505_),
    .B1(_0506_),
    .B2(\mod.registers.r2[3] ),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3685_ (.A1(\mod.registers.r4[3] ),
    .A2(_0508_),
    .B(_0421_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3686_ (.A1(_0652_),
    .A2(_0653_),
    .A3(_0654_),
    .A4(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3687_ (.A1(\mod.registers.r5[3] ),
    .A2(_0547_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3688_ (.A1(\mod.registers.r7[3] ),
    .A2(_0548_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3689_ (.A1(\mod.registers.r9[3] ),
    .A2(_0544_),
    .B1(_0545_),
    .B2(\mod.registers.r3[3] ),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3690_ (.I(\mod.registers.r12[3] ),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3691_ (.I(_0417_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3692_ (.I(\mod.registers.r15[3] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3693_ (.A1(_0660_),
    .A2(_0433_),
    .A3(_0661_),
    .B1(_0563_),
    .B2(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3694_ (.A1(\mod.registers.r13[3] ),
    .A2(_0541_),
    .B1(_0542_),
    .B2(\mod.registers.r1[3] ),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3695_ (.A1(_0657_),
    .A2(_0658_),
    .A3(_0659_),
    .A4(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3696_ (.A1(_0651_),
    .A2(_0464_),
    .B1(_0656_),
    .B2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3697_ (.A1(_0528_),
    .A2(_0552_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3698_ (.I0(_0650_),
    .I1(_0666_),
    .S(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3699_ (.I(\mod.pc_2[1] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3700_ (.A1(\mod.registers.r1[1] ),
    .A2(_0521_),
    .B1(_0412_),
    .B2(\mod.registers.r2[1] ),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3701_ (.A1(\mod.registers.r13[1] ),
    .A2(_0520_),
    .B1(_3272_),
    .B2(\mod.registers.r8[1] ),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3702_ (.A1(\mod.registers.r6[1] ),
    .A2(_0503_),
    .B1(_0515_),
    .B2(\mod.registers.r12[1] ),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3703_ (.A1(\mod.registers.r4[1] ),
    .A2(_0419_),
    .B(_3264_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3704_ (.A1(_0670_),
    .A2(_0671_),
    .A3(_0672_),
    .A4(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3705_ (.A1(\mod.registers.r15[1] ),
    .A2(_0514_),
    .B1(_0512_),
    .B2(\mod.registers.r3[1] ),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3706_ (.A1(\mod.registers.r14[1] ),
    .A2(_0502_),
    .B1(_3291_),
    .B2(\mod.registers.r11[1] ),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3707_ (.A1(\mod.registers.r5[1] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\mod.registers.r7[1] ),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3708_ (.A1(\mod.registers.r9[1] ),
    .A2(_0511_),
    .B1(_0500_),
    .B2(\mod.registers.r10[1] ),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3709_ (.A1(_0675_),
    .A2(_0676_),
    .A3(_0677_),
    .A4(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3710_ (.A1(_0669_),
    .A2(_0528_),
    .B1(_0674_),
    .B2(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3711_ (.I(_3261_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3712_ (.A1(_0579_),
    .A2(_0680_),
    .A3(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3713_ (.I(_0556_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3714_ (.I(_0557_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3715_ (.A1(_0683_),
    .A2(_0684_),
    .B(_0453_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3716_ (.A1(_0682_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3717_ (.I(_0615_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3718_ (.A1(_0687_),
    .A2(_0492_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3719_ (.A1(_0470_),
    .A2(_0488_),
    .B(_0560_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3720_ (.A1(_0688_),
    .A2(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3721_ (.I(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3722_ (.A1(_0691_),
    .A2(_0622_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3723_ (.A1(_0627_),
    .A2(_0668_),
    .B1(_0686_),
    .B2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3724_ (.I(_0471_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3725_ (.A1(\mod.registers.r3[3] ),
    .A2(_0694_),
    .B1(_0596_),
    .B2(\mod.registers.r7[3] ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3726_ (.I(_0465_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3727_ (.I(_0466_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3728_ (.A1(\mod.registers.r4[3] ),
    .A2(_0696_),
    .B1(_0697_),
    .B2(\mod.registers.r1[3] ),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(_0695_),
    .A2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3730_ (.I(_3185_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3731_ (.I(_3190_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3732_ (.A1(\mod.registers.r6[3] ),
    .A2(_0700_),
    .B1(_0468_),
    .B2(\mod.registers.r5[3] ),
    .C1(\mod.registers.r2[3] ),
    .C2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3733_ (.I(_3198_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3734_ (.A1(\mod.registers.r10[3] ),
    .A2(_0602_),
    .B1(_0703_),
    .B2(\mod.registers.r9[3] ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3735_ (.I(_3202_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3736_ (.I(_3204_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3737_ (.A1(\mod.registers.r11[3] ),
    .A2(_0705_),
    .B1(_0706_),
    .B2(\mod.registers.r8[3] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3738_ (.A1(_0660_),
    .A2(_3213_),
    .A3(_3214_),
    .B1(_3218_),
    .B2(_0662_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3739_ (.A1(\mod.registers.r14[3] ),
    .A2(_0607_),
    .B1(_0608_),
    .B2(\mod.registers.r13[3] ),
    .C(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3740_ (.A1(_0702_),
    .A2(_0704_),
    .A3(_0707_),
    .A4(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3741_ (.I(_3215_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3742_ (.I0(\mod.funct7[0] ),
    .I1(_0711_),
    .S(_0617_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3743_ (.A1(_0615_),
    .A2(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3744_ (.A1(_0595_),
    .A2(_0699_),
    .A3(_0710_),
    .B(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3745_ (.A1(_3246_),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3746_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3747_ (.I(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3748_ (.A1(_0624_),
    .A2(_0693_),
    .B(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3749_ (.A1(_0595_),
    .A2(_0699_),
    .A3(_0710_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3750_ (.I(_0560_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3751_ (.A1(_0720_),
    .A2(_0712_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3752_ (.A1(_3239_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3753_ (.A1(_0719_),
    .A2(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3754_ (.I(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3755_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3756_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3757_ (.I(\mod.pc_2[12] ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3758_ (.I(_3266_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3759_ (.I(_3272_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3760_ (.I(_0500_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3761_ (.A1(\mod.registers.r8[12] ),
    .A2(_0729_),
    .B1(_0730_),
    .B2(\mod.registers.r10[12] ),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3762_ (.I(_0502_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3763_ (.I(_0503_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3764_ (.A1(\mod.registers.r14[12] ),
    .A2(_0732_),
    .B1(_0733_),
    .B2(\mod.registers.r6[12] ),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3765_ (.I(_3291_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3766_ (.I(_0412_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3767_ (.A1(\mod.registers.r11[12] ),
    .A2(_0735_),
    .B1(_0736_),
    .B2(\mod.registers.r2[12] ),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3768_ (.I(_0419_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3769_ (.A1(\mod.registers.r4[12] ),
    .A2(_0738_),
    .B(_3266_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3770_ (.A1(_0731_),
    .A2(_0734_),
    .A3(_0737_),
    .A4(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3771_ (.I(_0517_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3772_ (.A1(\mod.registers.r5[12] ),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3773_ (.I(_0518_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3774_ (.A1(\mod.registers.r7[12] ),
    .A2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3775_ (.I(_0520_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3776_ (.I(_0521_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3777_ (.I(\mod.registers.r12[12] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3778_ (.I(\mod.registers.r15[12] ),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3779_ (.A1(_0747_),
    .A2(_0433_),
    .A3(_0661_),
    .B1(_0563_),
    .B2(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3780_ (.A1(\mod.registers.r13[12] ),
    .A2(_0745_),
    .B1(_0746_),
    .B2(\mod.registers.r1[12] ),
    .C(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3781_ (.I(_0511_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3782_ (.I(_0512_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3783_ (.A1(\mod.registers.r9[12] ),
    .A2(_0751_),
    .B1(_0752_),
    .B2(\mod.registers.r3[12] ),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3784_ (.A1(_0742_),
    .A2(_0744_),
    .A3(_0750_),
    .A4(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3785_ (.A1(_0727_),
    .A2(_0728_),
    .B1(_0740_),
    .B2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3786_ (.A1(_0683_),
    .A2(_0684_),
    .B(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3787_ (.I(_0728_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3788_ (.I(\mod.pc_2[13] ),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3789_ (.I(_0458_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3790_ (.A1(\mod.registers.r8[13] ),
    .A2(_3273_),
    .B1(_3279_),
    .B2(\mod.registers.r10[13] ),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3791_ (.A1(\mod.registers.r14[13] ),
    .A2(_3283_),
    .B1(_3287_),
    .B2(\mod.registers.r6[13] ),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3792_ (.A1(\mod.registers.r11[13] ),
    .A2(_0735_),
    .B1(_0736_),
    .B2(\mod.registers.r2[13] ),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3793_ (.A1(\mod.registers.r4[13] ),
    .A2(_0738_),
    .B(_3238_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3794_ (.A1(_0760_),
    .A2(_0761_),
    .A3(_0762_),
    .A4(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3795_ (.I(_0514_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3796_ (.I(_0515_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3797_ (.A1(\mod.registers.r15[13] ),
    .A2(_0765_),
    .B1(_0766_),
    .B2(\mod.registers.r12[13] ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3798_ (.A1(\mod.registers.r13[13] ),
    .A2(_0447_),
    .B1(_0449_),
    .B2(\mod.registers.r1[13] ),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3799_ (.A1(\mod.registers.r9[13] ),
    .A2(_0428_),
    .B1(_0752_),
    .B2(\mod.registers.r3[13] ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3800_ (.A1(\mod.registers.r5[13] ),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\mod.registers.r7[13] ),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3801_ (.A1(_0767_),
    .A2(_0768_),
    .A3(_0769_),
    .A4(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3802_ (.A1(_0758_),
    .A2(_0759_),
    .B1(_0764_),
    .B2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3803_ (.I(_0772_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3804_ (.I(_0552_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3805_ (.A1(_0757_),
    .A2(_0773_),
    .A3(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3806_ (.A1(_0756_),
    .A2(_0775_),
    .B(_0496_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3807_ (.I(_0498_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3808_ (.I(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3809_ (.I(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3810_ (.A1(\mod.registers.r5[14] ),
    .A2(_0741_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3811_ (.A1(\mod.registers.r15[14] ),
    .A2(_0765_),
    .B1(_0751_),
    .B2(\mod.registers.r9[14] ),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3812_ (.A1(\mod.registers.r3[14] ),
    .A2(_0752_),
    .B1(_0736_),
    .B2(\mod.registers.r2[14] ),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3813_ (.A1(\mod.registers.r7[14] ),
    .A2(_0743_),
    .B1(_0729_),
    .B2(\mod.registers.r8[14] ),
    .C1(\mod.registers.r12[14] ),
    .C2(_0766_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3814_ (.A1(_0780_),
    .A2(_0781_),
    .A3(_0782_),
    .A4(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3815_ (.A1(\mod.registers.r11[14] ),
    .A2(_0735_),
    .B1(_0746_),
    .B2(\mod.registers.r1[14] ),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3816_ (.A1(\mod.registers.r13[14] ),
    .A2(_0745_),
    .B1(_0738_),
    .B2(\mod.registers.r4[14] ),
    .C1(_0733_),
    .C2(\mod.registers.r6[14] ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3817_ (.A1(\mod.registers.r14[14] ),
    .A2(_0732_),
    .B1(_0730_),
    .B2(\mod.registers.r10[14] ),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3818_ (.A1(_0785_),
    .A2(_0786_),
    .A3(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3819_ (.A1(_0784_),
    .A2(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3820_ (.A1(_0779_),
    .A2(_0789_),
    .B1(_0556_),
    .B2(_0557_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3821_ (.A1(\mod.registers.r13[15] ),
    .A2(_0745_),
    .B1(_0732_),
    .B2(\mod.registers.r14[15] ),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3822_ (.A1(\mod.registers.r5[15] ),
    .A2(_0440_),
    .B1(_0442_),
    .B2(\mod.registers.r7[15] ),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3823_ (.A1(\mod.registers.r6[15] ),
    .A2(_0733_),
    .B1(_0766_),
    .B2(\mod.registers.r12[15] ),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3824_ (.A1(\mod.registers.r1[15] ),
    .A2(_0746_),
    .B1(_0431_),
    .B2(\mod.registers.r3[15] ),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3825_ (.A1(\mod.registers.r9[15] ),
    .A2(_0751_),
    .B1(_0730_),
    .B2(\mod.registers.r10[15] ),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3826_ (.A1(_0792_),
    .A2(_0793_),
    .A3(_0794_),
    .A4(_0795_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3827_ (.A1(\mod.registers.r11[15] ),
    .A2(_0735_),
    .B1(_0738_),
    .B2(\mod.registers.r4[15] ),
    .C1(_0736_),
    .C2(\mod.registers.r2[15] ),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3828_ (.A1(\mod.registers.r8[15] ),
    .A2(_0729_),
    .B1(_0765_),
    .B2(\mod.registers.r15[15] ),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3829_ (.A1(_0791_),
    .A2(_0796_),
    .A3(_0797_),
    .A4(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3830_ (.A1(_0579_),
    .A2(_0799_),
    .A3(_3262_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_0690_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3832_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3833_ (.A1(_0790_),
    .A2(_0800_),
    .B(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3834_ (.A1(_3253_),
    .A2(_0599_),
    .A3(_0613_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3835_ (.A1(_0560_),
    .A2(_0618_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3836_ (.A1(_0577_),
    .A2(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3837_ (.A1(_0804_),
    .A2(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3838_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3839_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3840_ (.A1(_0776_),
    .A2(_0803_),
    .B(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3841_ (.I(_0622_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3842_ (.I(_0801_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3843_ (.I(_0556_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3844_ (.I(_0557_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3845_ (.A1(\mod.registers.r8[11] ),
    .A2(_0531_),
    .B1(_0500_),
    .B2(\mod.registers.r10[11] ),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3846_ (.A1(\mod.registers.r14[11] ),
    .A2(_0502_),
    .B1(_0503_),
    .B2(\mod.registers.r6[11] ),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3847_ (.A1(\mod.registers.r11[11] ),
    .A2(_0505_),
    .B1(_0412_),
    .B2(\mod.registers.r2[11] ),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3848_ (.A1(\mod.registers.r4[11] ),
    .A2(_0419_),
    .B(_3264_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3849_ (.A1(_0815_),
    .A2(_0816_),
    .A3(_0817_),
    .A4(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3850_ (.A1(\mod.registers.r15[11] ),
    .A2(_0514_),
    .B1(_0515_),
    .B2(\mod.registers.r12[11] ),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3851_ (.A1(\mod.registers.r9[11] ),
    .A2(_0511_),
    .B1(_0512_),
    .B2(\mod.registers.r3[11] ),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3852_ (.A1(\mod.registers.r5[11] ),
    .A2(_0517_),
    .B1(_0518_),
    .B2(\mod.registers.r7[11] ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3853_ (.A1(\mod.registers.r13[11] ),
    .A2(_0520_),
    .B1(_0521_),
    .B2(\mod.registers.r1[11] ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3854_ (.A1(_0820_),
    .A2(_0821_),
    .A3(_0822_),
    .A4(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3855_ (.A1(\mod.pc_2[11] ),
    .A2(_0777_),
    .B1(_0819_),
    .B2(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3856_ (.I(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3857_ (.A1(_0813_),
    .A2(_0814_),
    .A3(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3858_ (.I(_0728_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3859_ (.A1(\mod.registers.r8[10] ),
    .A2(_0729_),
    .B1(_0730_),
    .B2(\mod.registers.r10[10] ),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3860_ (.A1(\mod.registers.r14[10] ),
    .A2(_0732_),
    .B1(_0733_),
    .B2(\mod.registers.r6[10] ),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3861_ (.A1(\mod.registers.r11[10] ),
    .A2(_3292_),
    .B1(_0413_),
    .B2(\mod.registers.r2[10] ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3862_ (.A1(\mod.registers.r4[10] ),
    .A2(_0420_),
    .B(_3265_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3863_ (.A1(_0829_),
    .A2(_0830_),
    .A3(_0831_),
    .A4(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3864_ (.A1(\mod.registers.r9[10] ),
    .A2(_0751_),
    .B1(_0752_),
    .B2(\mod.registers.r3[10] ),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3865_ (.A1(\mod.registers.r15[10] ),
    .A2(_0765_),
    .B1(_0766_),
    .B2(\mod.registers.r12[10] ),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3866_ (.A1(\mod.registers.r5[10] ),
    .A2(_0741_),
    .B1(_0743_),
    .B2(\mod.registers.r7[10] ),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3867_ (.A1(\mod.registers.r13[10] ),
    .A2(_0745_),
    .B1(_0746_),
    .B2(\mod.registers.r1[10] ),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3868_ (.A1(_0834_),
    .A2(_0835_),
    .A3(_0836_),
    .A4(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3869_ (.A1(\mod.pc_2[10] ),
    .A2(_0778_),
    .B1(_0833_),
    .B2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3870_ (.I(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3871_ (.A1(_0828_),
    .A2(_0553_),
    .B(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3872_ (.A1(_0812_),
    .A2(_0827_),
    .A3(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3873_ (.I(\mod.pc_2[8] ),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3874_ (.A1(\mod.registers.r4[8] ),
    .A2(_0420_),
    .B1(_0435_),
    .B2(\mod.registers.r15[8] ),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3875_ (.A1(\mod.registers.r7[8] ),
    .A2(_0442_),
    .B1(_3287_),
    .B2(\mod.registers.r6[8] ),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3876_ (.I(_0631_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3877_ (.A1(_0846_),
    .A2(_0632_),
    .A3(\mod.registers.r11[8] ),
    .A4(_0634_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3878_ (.A1(_0631_),
    .A2(_0562_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3879_ (.A1(\mod.registers.r12[8] ),
    .A2(_0848_),
    .A3(_0638_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3880_ (.A1(_0846_),
    .A2(_0632_),
    .A3(\mod.registers.r8[8] ),
    .A4(_0638_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3881_ (.A1(_0777_),
    .A2(_0847_),
    .A3(_0849_),
    .A4(_0850_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3882_ (.A1(_0844_),
    .A2(_0845_),
    .A3(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3883_ (.A1(\mod.registers.r1[8] ),
    .A2(_0449_),
    .B1(_0431_),
    .B2(\mod.registers.r3[8] ),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3884_ (.A1(\mod.registers.r13[8] ),
    .A2(_0447_),
    .B1(_3279_),
    .B2(\mod.registers.r10[8] ),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3885_ (.A1(\mod.registers.r14[8] ),
    .A2(_3283_),
    .B1(_0428_),
    .B2(\mod.registers.r9[8] ),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3886_ (.A1(\mod.registers.r5[8] ),
    .A2(_0440_),
    .B1(_0413_),
    .B2(\mod.registers.r2[8] ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3887_ (.A1(_0853_),
    .A2(_0854_),
    .A3(_0855_),
    .A4(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3888_ (.A1(_0843_),
    .A2(_3239_),
    .B1(_0852_),
    .B2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3889_ (.I(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3890_ (.A1(_0813_),
    .A2(_0814_),
    .B(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3891_ (.I(_0552_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3892_ (.I(\mod.pc_2[9] ),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3893_ (.A1(\mod.registers.r8[9] ),
    .A2(_3273_),
    .B1(_0532_),
    .B2(\mod.registers.r10[9] ),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3894_ (.A1(\mod.registers.r14[9] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\mod.registers.r6[9] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3895_ (.A1(\mod.registers.r11[9] ),
    .A2(_3292_),
    .B1(_0506_),
    .B2(\mod.registers.r2[9] ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3896_ (.A1(\mod.registers.r4[9] ),
    .A2(_0508_),
    .B(_0421_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3897_ (.A1(_0863_),
    .A2(_0864_),
    .A3(_0865_),
    .A4(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3898_ (.A1(\mod.registers.r15[9] ),
    .A2(_0435_),
    .B1(_0437_),
    .B2(\mod.registers.r12[9] ),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3899_ (.A1(\mod.registers.r13[9] ),
    .A2(_0541_),
    .B1(_0542_),
    .B2(\mod.registers.r1[9] ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3900_ (.A1(\mod.registers.r9[9] ),
    .A2(_0544_),
    .B1(_0545_),
    .B2(\mod.registers.r3[9] ),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3901_ (.A1(\mod.registers.r5[9] ),
    .A2(_0547_),
    .B1(_0548_),
    .B2(\mod.registers.r7[9] ),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3902_ (.A1(_0868_),
    .A2(_0869_),
    .A3(_0870_),
    .A4(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3903_ (.A1(_0862_),
    .A2(_0464_),
    .B1(_0867_),
    .B2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3904_ (.I(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3905_ (.A1(_0828_),
    .A2(_0861_),
    .A3(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3906_ (.A1(_0802_),
    .A2(_0860_),
    .A3(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3907_ (.A1(_0811_),
    .A2(_0842_),
    .A3(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3908_ (.I(_0799_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3909_ (.I(_3170_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3910_ (.A1(\mod.registers.r7[4] ),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3911_ (.A1(\mod.registers.r3[4] ),
    .A2(_3165_),
    .B1(_0697_),
    .B2(\mod.registers.r1[4] ),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3912_ (.I(_3188_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3913_ (.A1(\mod.registers.r5[4] ),
    .A2(_0882_),
    .B1(_0706_),
    .B2(\mod.registers.r8[4] ),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3914_ (.I(_0485_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _3915_ (.A1(\mod.registers.r15[4] ),
    .A2(_0884_),
    .B1(_0600_),
    .B2(\mod.registers.r6[4] ),
    .C1(_0603_),
    .C2(\mod.registers.r9[4] ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3916_ (.A1(_0880_),
    .A2(_0881_),
    .A3(_0883_),
    .A4(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3917_ (.A1(_3172_),
    .A2(_3214_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3918_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3919_ (.I(_3211_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3920_ (.A1(\mod.registers.r12[4] ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\mod.registers.r13[4] ),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3921_ (.I(_3208_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3922_ (.A1(\mod.registers.r14[4] ),
    .A2(_0891_),
    .B1(_0705_),
    .B2(\mod.registers.r11[4] ),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3923_ (.I(_3191_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3924_ (.A1(\mod.registers.r2[4] ),
    .A2(_0893_),
    .B1(_3174_),
    .B2(\mod.registers.r4[4] ),
    .C1(\mod.registers.r10[4] ),
    .C2(_0602_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3925_ (.A1(_0890_),
    .A2(_0892_),
    .A3(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3926_ (.A1(_3253_),
    .A2(_0886_),
    .A3(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3927_ (.I0(\mod.funct7[1] ),
    .I1(\mod.funct7[0] ),
    .S(_0617_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3928_ (.A1(_0720_),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3929_ (.A1(_0759_),
    .A2(_0896_),
    .A3(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3930_ (.A1(_0878_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3931_ (.I(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3932_ (.I(_0457_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3933_ (.I(_3230_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3934_ (.I(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(_3231_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3936_ (.I(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3937_ (.A1(_0904_),
    .A2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3938_ (.A1(_0902_),
    .A2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3939_ (.A1(\mod.funct7[1] ),
    .A2(_0905_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3940_ (.A1(_3227_),
    .A2(_0902_),
    .B(_0909_),
    .C(_0903_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3941_ (.A1(_0908_),
    .A2(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3942_ (.I(_0911_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3943_ (.A1(_0726_),
    .A2(_0810_),
    .A3(_0877_),
    .B1(_0901_),
    .B2(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3944_ (.I(\mod.funct3[0] ),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3945_ (.A1(_3228_),
    .A2(_3233_),
    .A3(_0728_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3946_ (.A1(_0914_),
    .A2(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3947_ (.A1(_3227_),
    .A2(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3948_ (.I(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3949_ (.A1(_0718_),
    .A2(_0913_),
    .B(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3950_ (.A1(_3248_),
    .A2(_0916_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3951_ (.A1(_0724_),
    .A2(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3952_ (.I(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3953_ (.I(_0625_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3954_ (.A1(_0923_),
    .A2(_0808_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3955_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_3246_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3957_ (.A1(_0926_),
    .A2(_0774_),
    .B(_0453_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3958_ (.A1(_0925_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3959_ (.A1(_0455_),
    .A2(_0459_),
    .A3(_0452_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3960_ (.A1(_3248_),
    .A2(_0914_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3961_ (.A1(_3228_),
    .A2(_3240_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3962_ (.I(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3963_ (.A1(_0930_),
    .A2(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3964_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3965_ (.I(\mod.funct3[0] ),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3966_ (.A1(_3226_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3967_ (.A1(_0931_),
    .A2(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3968_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3969_ (.A1(_3233_),
    .A2(_0926_),
    .A3(_3249_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3970_ (.I(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3971_ (.A1(_0929_),
    .A2(_0934_),
    .B1(_0685_),
    .B2(_0938_),
    .C(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3972_ (.I(_3248_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3973_ (.I(_0935_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3974_ (.A1(_0942_),
    .A2(_0943_),
    .A3(_0915_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3975_ (.I(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3976_ (.A1(_3241_),
    .A2(_0945_),
    .B(_0463_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3977_ (.A1(_0922_),
    .A2(_0928_),
    .B(_0941_),
    .C(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3978_ (.A1(_3250_),
    .A2(_0463_),
    .B1(_0919_),
    .B2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3979_ (.A1(_3243_),
    .A2(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_0779_),
    .A2(_0878_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3981_ (.I(_3196_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3982_ (.A1(_3232_),
    .A2(_3252_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3983_ (.I(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3984_ (.I(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3985_ (.I(\mod.funct7[2] ),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3986_ (.A1(_0955_),
    .A2(_0952_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3987_ (.I(_0956_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3988_ (.A1(_0951_),
    .A2(_0954_),
    .B(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3989_ (.I(_3165_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3990_ (.I(_0701_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3991_ (.A1(\mod.registers.r3[15] ),
    .A2(_0959_),
    .B1(_0960_),
    .B2(\mod.registers.r2[15] ),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3992_ (.I(_0888_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3993_ (.I(_0485_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3994_ (.I(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3995_ (.A1(\mod.registers.r12[15] ),
    .A2(_0962_),
    .B1(_0964_),
    .B2(\mod.registers.r15[15] ),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3996_ (.I(_0600_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3997_ (.I(_0468_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3998_ (.I(_0473_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3999_ (.A1(\mod.registers.r6[15] ),
    .A2(_0966_),
    .B1(_0967_),
    .B2(\mod.registers.r5[15] ),
    .C1(_0968_),
    .C2(\mod.registers.r8[15] ),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4000_ (.A1(_0961_),
    .A2(_0965_),
    .A3(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4001_ (.I(_3174_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4002_ (.I(_0602_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4003_ (.A1(\mod.registers.r4[15] ),
    .A2(_0971_),
    .B1(_0972_),
    .B2(\mod.registers.r10[15] ),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4004_ (.I(_0605_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4005_ (.I(_3178_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4006_ (.A1(\mod.registers.r11[15] ),
    .A2(_0974_),
    .B1(_0975_),
    .B2(\mod.registers.r1[15] ),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4007_ (.I(_0607_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4008_ (.I(_3170_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4009_ (.A1(\mod.registers.r14[15] ),
    .A2(_0977_),
    .B1(_0978_),
    .B2(\mod.registers.r7[15] ),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4010_ (.I(_0608_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4011_ (.I(_0603_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4012_ (.A1(\mod.registers.r13[15] ),
    .A2(_0980_),
    .B1(_0981_),
    .B2(\mod.registers.r9[15] ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4013_ (.A1(_0973_),
    .A2(_0976_),
    .A3(_0979_),
    .A4(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4014_ (.A1(_0970_),
    .A2(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4015_ (.A1(_0955_),
    .A2(_0561_),
    .B(_0720_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4016_ (.A1(_0687_),
    .A2(_0984_),
    .B(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4017_ (.A1(_3247_),
    .A2(_0958_),
    .B(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4018_ (.A1(_0950_),
    .A2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4019_ (.I(_0799_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4020_ (.A1(_0989_),
    .A2(_0986_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4021_ (.A1(_0988_),
    .A2(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4022_ (.I(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4023_ (.A1(\mod.registers.r4[14] ),
    .A2(_0971_),
    .B1(_0975_),
    .B2(\mod.registers.r1[14] ),
    .C1(_0972_),
    .C2(\mod.registers.r10[14] ),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4024_ (.A1(\mod.registers.r14[14] ),
    .A2(_0977_),
    .B1(_0978_),
    .B2(\mod.registers.r7[14] ),
    .C1(_0981_),
    .C2(\mod.registers.r9[14] ),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4025_ (.A1(\mod.registers.r11[14] ),
    .A2(_0974_),
    .B1(_0980_),
    .B2(\mod.registers.r13[14] ),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4026_ (.A1(_0993_),
    .A2(_0994_),
    .A3(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4027_ (.A1(\mod.registers.r6[14] ),
    .A2(_0966_),
    .B1(_0967_),
    .B2(\mod.registers.r5[14] ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4028_ (.A1(\mod.registers.r15[14] ),
    .A2(_0964_),
    .B1(_0968_),
    .B2(\mod.registers.r8[14] ),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4029_ (.A1(\mod.registers.r3[14] ),
    .A2(_0959_),
    .B1(_0960_),
    .B2(\mod.registers.r2[14] ),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4030_ (.A1(_0997_),
    .A2(_0998_),
    .A3(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4031_ (.A1(\mod.registers.r12[14] ),
    .A2(_0962_),
    .B(_0996_),
    .C(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4032_ (.A1(\mod.funct7[2] ),
    .A2(_0614_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4033_ (.A1(_0687_),
    .A2(_1001_),
    .B(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4034_ (.A1(_0779_),
    .A2(_1003_),
    .A3(_0789_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4035_ (.A1(\mod.registers.r15[7] ),
    .A2(_0963_),
    .B1(_3186_),
    .B2(\mod.registers.r6[7] ),
    .C1(_3189_),
    .C2(\mod.registers.r5[7] ),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4036_ (.A1(\mod.registers.r2[7] ),
    .A2(_0701_),
    .B1(_3195_),
    .B2(\mod.registers.r10[7] ),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4037_ (.A1(\mod.registers.r11[7] ),
    .A2(_0605_),
    .B1(_3199_),
    .B2(\mod.registers.r9[7] ),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4038_ (.A1(_1005_),
    .A2(_1006_),
    .A3(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4039_ (.A1(\mod.registers.r12[7] ),
    .A2(_0888_),
    .B1(_0608_),
    .B2(\mod.registers.r13[7] ),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4040_ (.I(_0476_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4041_ (.A1(_3215_),
    .A2(_3168_),
    .A3(\mod.registers.r8[7] ),
    .A4(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4042_ (.A1(_0951_),
    .A2(_3216_),
    .A3(\mod.registers.r4[7] ),
    .A4(_1010_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4043_ (.A1(_3209_),
    .A2(_3217_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4044_ (.A1(_3166_),
    .A2(_3216_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4045_ (.I(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4046_ (.A1(\mod.registers.r3[7] ),
    .A2(_1013_),
    .A3(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4047_ (.A1(_0482_),
    .A2(_0483_),
    .A3(\mod.registers.r1[7] ),
    .A4(_1014_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4048_ (.A1(_1011_),
    .A2(_1012_),
    .A3(_1016_),
    .A4(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4049_ (.A1(\mod.registers.r14[7] ),
    .A2(_0607_),
    .B1(_0596_),
    .B2(\mod.registers.r7[7] ),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4050_ (.A1(_1009_),
    .A2(_1018_),
    .A3(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4051_ (.A1(_3264_),
    .A2(_1002_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4052_ (.A1(_3254_),
    .A2(_1008_),
    .A3(_1020_),
    .B(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4053_ (.A1(_3232_),
    .A2(_3251_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4054_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4055_ (.I0(_3226_),
    .I1(_0618_),
    .S(_1024_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4056_ (.A1(_0458_),
    .A2(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4057_ (.A1(_0533_),
    .A2(_0536_),
    .A3(_0537_),
    .A4(_0538_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4058_ (.A1(_0540_),
    .A2(_0543_),
    .A3(_0546_),
    .A4(_0549_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4059_ (.A1(\mod.pc_2[7] ),
    .A2(_0499_),
    .B1(_1027_),
    .B2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4060_ (.A1(_1022_),
    .A2(_1026_),
    .B(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4061_ (.A1(_1029_),
    .A2(_1022_),
    .A3(_1026_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4062_ (.A1(_1030_),
    .A2(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4063_ (.I(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4064_ (.A1(\mod.registers.r11[6] ),
    .A2(_3202_),
    .B1(_3194_),
    .B2(\mod.registers.r10[6] ),
    .C1(\mod.registers.r2[6] ),
    .C2(_3190_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4065_ (.A1(\mod.registers.r15[6] ),
    .A2(_0963_),
    .B1(_3186_),
    .B2(\mod.registers.r6[6] ),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4066_ (.A1(\mod.registers.r5[6] ),
    .A2(_3189_),
    .B1(_3199_),
    .B2(\mod.registers.r9[6] ),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4067_ (.A1(_1034_),
    .A2(_1035_),
    .A3(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4068_ (.A1(\mod.registers.r3[6] ),
    .A2(_0471_),
    .B1(_0465_),
    .B2(\mod.registers.r4[6] ),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4069_ (.A1(\mod.registers.r1[6] ),
    .A2(_0466_),
    .B1(_3204_),
    .B2(\mod.registers.r8[6] ),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4070_ (.A1(\mod.registers.r14[6] ),
    .A2(_3208_),
    .B1(_3169_),
    .B2(\mod.registers.r7[6] ),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4071_ (.A1(\mod.registers.r12[6] ),
    .A2(_0887_),
    .B1(_3211_),
    .B2(\mod.registers.r13[6] ),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4072_ (.A1(_1038_),
    .A2(_1039_),
    .A3(_1040_),
    .A4(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4073_ (.A1(_0489_),
    .A2(_1037_),
    .A3(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4074_ (.I(_1024_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4075_ (.A1(\mod.funct3[1] ),
    .A2(_1024_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4076_ (.A1(_1044_),
    .A2(_0491_),
    .B(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4077_ (.A1(_1021_),
    .A2(_1043_),
    .B1(_1046_),
    .B2(_0458_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4078_ (.A1(_0524_),
    .A2(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4079_ (.I(_1048_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4080_ (.A1(_1033_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4081_ (.I(\mod.pc_2[2] ),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4082_ (.A1(_0629_),
    .A2(_0630_),
    .A3(_0642_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4083_ (.A1(_0644_),
    .A2(_0645_),
    .A3(_0646_),
    .A4(_0648_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4084_ (.A1(_1051_),
    .A2(_0499_),
    .B1(_1052_),
    .B2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4085_ (.A1(_0759_),
    .A2(_0620_),
    .A3(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4086_ (.I(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4087_ (.A1(_0652_),
    .A2(_0653_),
    .A3(_0654_),
    .A4(_0655_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4088_ (.A1(_0657_),
    .A2(_0658_),
    .A3(_0659_),
    .A4(_0664_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4089_ (.A1(\mod.pc_2[3] ),
    .A2(_0778_),
    .B1(_1057_),
    .B2(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4090_ (.A1(_0723_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4091_ (.A1(_0804_),
    .A2(_0806_),
    .B(_0650_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4092_ (.A1(_3245_),
    .A2(_0714_),
    .A3(_1059_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4093_ (.A1(_0719_),
    .A2(_0722_),
    .B(_0666_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4094_ (.A1(_1055_),
    .A2(_1061_),
    .A3(_1062_),
    .A4(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4095_ (.A1(_0670_),
    .A2(_0671_),
    .A3(_0672_),
    .A4(_0673_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4096_ (.A1(_0675_),
    .A2(_0676_),
    .A3(_0677_),
    .A4(_0678_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4097_ (.A1(\mod.pc_2[1] ),
    .A2(_0777_),
    .B1(_1065_),
    .B2(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4098_ (.A1(_0759_),
    .A2(_0494_),
    .A3(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4099_ (.I(_1067_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4100_ (.A1(_0688_),
    .A2(_0689_),
    .A3(_1069_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4101_ (.A1(_1068_),
    .A2(_0929_),
    .B(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4102_ (.I(_1062_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4103_ (.A1(_1056_),
    .A2(_1060_),
    .B1(_1064_),
    .B2(_1071_),
    .C(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4104_ (.A1(_0567_),
    .A2(_0572_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _4105_ (.A1(_0578_),
    .A2(_1074_),
    .A3(_0896_),
    .A4(_0898_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4106_ (.I(_0591_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4107_ (.A1(\mod.funct3[0] ),
    .A2(_1023_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4108_ (.A1(_1024_),
    .A2(_3259_),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4109_ (.A1(\mod.registers.r2[5] ),
    .A2(_3190_),
    .B1(_3169_),
    .B2(\mod.registers.r7[5] ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4110_ (.A1(\mod.registers.r3[5] ),
    .A2(_0471_),
    .B1(_0466_),
    .B2(\mod.registers.r1[5] ),
    .C1(_3201_),
    .C2(\mod.registers.r11[5] ),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4111_ (.A1(\mod.registers.r5[5] ),
    .A2(_3188_),
    .B1(_3211_),
    .B2(\mod.registers.r13[5] ),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4112_ (.A1(_1079_),
    .A2(_1080_),
    .A3(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4113_ (.A1(\mod.registers.r12[5] ),
    .A2(_0887_),
    .B1(_3185_),
    .B2(\mod.registers.r6[5] ),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4114_ (.A1(\mod.registers.r4[5] ),
    .A2(_0465_),
    .B1(_3194_),
    .B2(\mod.registers.r10[5] ),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4115_ (.A1(\mod.registers.r8[5] ),
    .A2(_3204_),
    .B1(_3198_),
    .B2(\mod.registers.r9[5] ),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4116_ (.A1(\mod.registers.r15[5] ),
    .A2(_0485_),
    .B1(_3208_),
    .B2(\mod.registers.r14[5] ),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4117_ (.A1(_1083_),
    .A2(_1084_),
    .A3(_1085_),
    .A4(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4118_ (.A1(_1082_),
    .A2(_1087_),
    .B(_0457_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4119_ (.I(\mod.funct7[2] ),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4120_ (.I(\mod.funct7[1] ),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4121_ (.I0(_1089_),
    .I1(_1090_),
    .S(_0617_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4122_ (.A1(_0615_),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4123_ (.A1(_3238_),
    .A2(_1078_),
    .B(_1088_),
    .C(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4124_ (.A1(_1076_),
    .A2(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4125_ (.A1(_0899_),
    .A2(_0574_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4126_ (.A1(_1075_),
    .A2(_1094_),
    .A3(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4127_ (.I(_1032_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4128_ (.A1(_1076_),
    .A2(_1093_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4129_ (.I(_1093_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4130_ (.A1(_1076_),
    .A2(_1099_),
    .B(_1075_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4131_ (.A1(_1097_),
    .A2(_1049_),
    .A3(_1098_),
    .A4(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4132_ (.A1(_1050_),
    .A2(_1073_),
    .A3(_1096_),
    .B(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4133_ (.I(_1047_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4134_ (.I(_1030_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4135_ (.A1(_1031_),
    .A2(_0525_),
    .A3(_1103_),
    .B(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4136_ (.I(_3195_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4137_ (.A1(\mod.registers.r10[9] ),
    .A2(_1106_),
    .B1(_0703_),
    .B2(\mod.registers.r9[9] ),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4138_ (.A1(\mod.registers.r3[9] ),
    .A2(_0694_),
    .B1(_0882_),
    .B2(\mod.registers.r5[9] ),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4139_ (.A1(_1107_),
    .A2(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4140_ (.I(_0888_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(\mod.registers.r12[9] ),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4142_ (.A1(\mod.registers.r2[9] ),
    .A2(_0701_),
    .B1(_3178_),
    .B2(\mod.registers.r1[9] ),
    .C1(_0596_),
    .C2(\mod.registers.r7[9] ),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4143_ (.I(_3168_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4144_ (.A1(_3215_),
    .A2(_1113_),
    .A3(\mod.registers.r11[9] ),
    .A4(_1013_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4145_ (.A1(_0480_),
    .A2(_3256_),
    .A3(\mod.registers.r14[9] ),
    .A4(_0478_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4146_ (.A1(_0482_),
    .A2(_0483_),
    .A3(\mod.registers.r13[9] ),
    .A4(_0478_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4147_ (.A1(_0951_),
    .A2(_0616_),
    .A3(\mod.registers.r4[9] ),
    .A4(_1010_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4148_ (.A1(_1114_),
    .A2(_1115_),
    .A3(_1116_),
    .A4(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4149_ (.A1(\mod.registers.r15[9] ),
    .A2(_0884_),
    .B1(_0600_),
    .B2(\mod.registers.r6[9] ),
    .C1(_0473_),
    .C2(\mod.registers.r8[9] ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4150_ (.A1(_1111_),
    .A2(_1112_),
    .A3(_1118_),
    .A4(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4151_ (.A1(_3253_),
    .A2(_1109_),
    .A3(_1120_),
    .B(_1021_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4152_ (.I0(_0637_),
    .I1(_0897_),
    .S(_1044_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4153_ (.A1(_0577_),
    .A2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4154_ (.A1(_1121_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_0873_),
    .A2(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4156_ (.A1(_0873_),
    .A2(_1124_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4157_ (.A1(_1125_),
    .A2(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4158_ (.I(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4159_ (.A1(\mod.registers.r12[8] ),
    .A2(_1110_),
    .B1(_0879_),
    .B2(\mod.registers.r7[8] ),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4160_ (.A1(\mod.registers.r14[8] ),
    .A2(_0891_),
    .B1(_0889_),
    .B2(\mod.registers.r13[8] ),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4161_ (.A1(_1129_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4162_ (.A1(\mod.registers.r10[8] ),
    .A2(_1106_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4163_ (.A1(\mod.registers.r6[8] ),
    .A2(_0700_),
    .B1(_0696_),
    .B2(\mod.registers.r4[8] ),
    .C1(_0603_),
    .C2(\mod.registers.r9[8] ),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4164_ (.A1(_0711_),
    .A2(_1113_),
    .A3(\mod.registers.r8[8] ),
    .A4(_1010_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4165_ (.I(_3183_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4166_ (.I(_0483_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4167_ (.A1(_1135_),
    .A2(_1136_),
    .A3(\mod.registers.r1[8] ),
    .A4(_1015_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4168_ (.A1(\mod.registers.r15[8] ),
    .A2(_0963_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4169_ (.A1(\mod.registers.r3[8] ),
    .A2(_1013_),
    .A3(_1015_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4170_ (.A1(_1134_),
    .A2(_1137_),
    .A3(_1138_),
    .A4(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4171_ (.A1(\mod.registers.r2[8] ),
    .A2(_0893_),
    .B1(_0468_),
    .B2(\mod.registers.r5[8] ),
    .C1(\mod.registers.r11[8] ),
    .C2(_0605_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4172_ (.A1(_1132_),
    .A2(_1133_),
    .A3(_1140_),
    .A4(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4173_ (.I(_1021_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4174_ (.A1(_0595_),
    .A2(_1131_),
    .A3(_1142_),
    .B(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4175_ (.I0(_0633_),
    .I1(_0712_),
    .S(_1044_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4176_ (.A1(_3266_),
    .A2(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(_1144_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4178_ (.A1(_0858_),
    .A2(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4179_ (.A1(_0858_),
    .A2(_1147_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4180_ (.A1(_1148_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4181_ (.I(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4182_ (.I(_0489_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4183_ (.A1(\mod.registers.r15[10] ),
    .A2(_0884_),
    .B1(_0879_),
    .B2(\mod.registers.r7[10] ),
    .C1(\mod.registers.r3[10] ),
    .C2(_0694_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4184_ (.A1(\mod.registers.r5[10] ),
    .A2(_0882_),
    .B1(_0696_),
    .B2(\mod.registers.r4[10] ),
    .C1(_0706_),
    .C2(\mod.registers.r8[10] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4185_ (.A1(\mod.registers.r12[10] ),
    .A2(_1110_),
    .B1(_1106_),
    .B2(\mod.registers.r10[10] ),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4186_ (.A1(_1153_),
    .A2(_1154_),
    .A3(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4187_ (.A1(\mod.registers.r1[10] ),
    .A2(_0697_),
    .B1(_0980_),
    .B2(\mod.registers.r13[10] ),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4188_ (.A1(\mod.registers.r6[10] ),
    .A2(_0700_),
    .B1(_0705_),
    .B2(\mod.registers.r11[10] ),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4189_ (.A1(\mod.registers.r14[10] ),
    .A2(_0891_),
    .B1(_0703_),
    .B2(\mod.registers.r9[10] ),
    .C1(\mod.registers.r2[10] ),
    .C2(_0893_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4190_ (.A1(_1157_),
    .A2(_1158_),
    .A3(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4191_ (.A1(_1152_),
    .A2(_1156_),
    .A3(_1160_),
    .B(_1143_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4192_ (.A1(_0636_),
    .A2(_0952_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4193_ (.A1(_0953_),
    .A2(_1091_),
    .B(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4194_ (.A1(_3245_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4195_ (.A1(_0839_),
    .A2(_1161_),
    .A3(_1164_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4196_ (.A1(_1161_),
    .A2(_1164_),
    .B(_0839_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4197_ (.A1(_1165_),
    .A2(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4198_ (.A1(\mod.registers.r14[11] ),
    .A2(_0891_),
    .B1(_0703_),
    .B2(\mod.registers.r9[11] ),
    .C1(\mod.registers.r2[11] ),
    .C2(_0893_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4199_ (.A1(\mod.registers.r11[11] ),
    .A2(_0705_),
    .B1(_0697_),
    .B2(\mod.registers.r1[11] ),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4200_ (.A1(\mod.registers.r6[11] ),
    .A2(_0700_),
    .B1(_0889_),
    .B2(\mod.registers.r13[11] ),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4201_ (.A1(_1168_),
    .A2(_1169_),
    .A3(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4202_ (.A1(\mod.registers.r3[11] ),
    .A2(_0694_),
    .B1(_0879_),
    .B2(\mod.registers.r7[11] ),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4203_ (.A1(\mod.registers.r15[11] ),
    .A2(_0884_),
    .B1(_1106_),
    .B2(\mod.registers.r10[11] ),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4204_ (.A1(\mod.registers.r8[11] ),
    .A2(_0706_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4205_ (.A1(\mod.registers.r12[11] ),
    .A2(_1110_),
    .B1(_0882_),
    .B2(\mod.registers.r5[11] ),
    .C1(_0696_),
    .C2(\mod.registers.r4[11] ),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4206_ (.A1(_1172_),
    .A2(_1173_),
    .A3(_1174_),
    .A4(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4207_ (.A1(_1152_),
    .A2(_1171_),
    .A3(_1176_),
    .B(_1143_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4208_ (.A1(_0424_),
    .A2(_0953_),
    .B(_0956_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4209_ (.A1(_3239_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4210_ (.A1(_1177_),
    .A2(_1179_),
    .B(_0826_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4211_ (.A1(_0825_),
    .A2(_1177_),
    .A3(_1179_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4212_ (.A1(_1180_),
    .A2(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4213_ (.A1(_1128_),
    .A2(_1151_),
    .A3(_1167_),
    .A4(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4214_ (.A1(_1102_),
    .A2(_1105_),
    .B(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4215_ (.I(_1166_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4216_ (.A1(_0874_),
    .A2(_1124_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4217_ (.A1(_0859_),
    .A2(_1147_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4218_ (.A1(_1186_),
    .A2(_1187_),
    .B(_1126_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4219_ (.A1(_1185_),
    .A2(_1188_),
    .B(_1181_),
    .C(_1165_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4220_ (.A1(_1180_),
    .A2(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4221_ (.I(_0720_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4222_ (.A1(\mod.registers.r15[13] ),
    .A2(_0964_),
    .B1(_0968_),
    .B2(\mod.registers.r8[13] ),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4223_ (.A1(\mod.registers.r6[13] ),
    .A2(_0966_),
    .B1(_0967_),
    .B2(\mod.registers.r5[13] ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4224_ (.A1(\mod.registers.r14[13] ),
    .A2(_0977_),
    .B1(_0889_),
    .B2(\mod.registers.r13[13] ),
    .C1(_0978_),
    .C2(\mod.registers.r7[13] ),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4225_ (.A1(\mod.registers.r1[13] ),
    .A2(_0975_),
    .B1(_0981_),
    .B2(\mod.registers.r9[13] ),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4226_ (.A1(_1192_),
    .A2(_1193_),
    .A3(_1194_),
    .A4(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4227_ (.A1(\mod.registers.r12[13] ),
    .A2(_0962_),
    .B1(_0959_),
    .B2(\mod.registers.r3[13] ),
    .C1(_0960_),
    .C2(\mod.registers.r2[13] ),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4228_ (.A1(\mod.registers.r11[13] ),
    .A2(_0974_),
    .B1(_0972_),
    .B2(\mod.registers.r10[13] ),
    .C1(\mod.registers.r4[13] ),
    .C2(_0971_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4229_ (.A1(_1197_),
    .A2(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4230_ (.A1(_1152_),
    .A2(_1196_),
    .A3(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4231_ (.A1(_1135_),
    .A2(_1191_),
    .A3(_0561_),
    .B1(_0985_),
    .B2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4232_ (.I(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4233_ (.A1(_0772_),
    .A2(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4234_ (.I(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4235_ (.I(_0778_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4236_ (.I(_1044_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4237_ (.I(_0956_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4238_ (.A1(_1136_),
    .A2(_1206_),
    .B(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4239_ (.A1(\mod.registers.r4[12] ),
    .A2(_0971_),
    .B1(_0972_),
    .B2(\mod.registers.r10[12] ),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4240_ (.A1(\mod.registers.r11[12] ),
    .A2(_0974_),
    .B1(_0980_),
    .B2(\mod.registers.r13[12] ),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4241_ (.A1(\mod.registers.r14[12] ),
    .A2(_0977_),
    .B1(_0978_),
    .B2(\mod.registers.r7[12] ),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4242_ (.A1(\mod.registers.r12[12] ),
    .A2(_0962_),
    .B1(_0975_),
    .B2(\mod.registers.r1[12] ),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4243_ (.A1(_1209_),
    .A2(_1210_),
    .A3(_1211_),
    .A4(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4244_ (.A1(\mod.registers.r3[12] ),
    .A2(_0959_),
    .B1(_0960_),
    .B2(\mod.registers.r2[12] ),
    .C1(_0964_),
    .C2(\mod.registers.r15[12] ),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4245_ (.A1(\mod.registers.r6[12] ),
    .A2(_0966_),
    .B1(_0967_),
    .B2(\mod.registers.r5[12] ),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4246_ (.A1(\mod.registers.r8[12] ),
    .A2(_0968_),
    .B1(_0981_),
    .B2(\mod.registers.r9[12] ),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4247_ (.A1(_1214_),
    .A2(_1215_),
    .A3(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4248_ (.A1(_1213_),
    .A2(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4249_ (.A1(_1152_),
    .A2(_1218_),
    .B(_1143_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4250_ (.A1(_1205_),
    .A2(_1208_),
    .B(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4251_ (.A1(_0755_),
    .A2(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4252_ (.A1(_0755_),
    .A2(_1220_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4253_ (.A1(_1221_),
    .A2(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4254_ (.I(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4255_ (.A1(_1184_),
    .A2(_1190_),
    .B(_1204_),
    .C(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4256_ (.I(_0773_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4257_ (.A1(_1226_),
    .A2(_1201_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4258_ (.I(_1221_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4259_ (.A1(_1226_),
    .A2(_1201_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4260_ (.A1(_1227_),
    .A2(_1228_),
    .B(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4261_ (.I(_1003_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4262_ (.A1(_0779_),
    .A2(_0789_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4263_ (.A1(_1113_),
    .A2(_0953_),
    .B(_0957_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4264_ (.A1(_0926_),
    .A2(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4265_ (.A1(_3247_),
    .A2(_1231_),
    .B(_1232_),
    .C(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4266_ (.A1(_1004_),
    .A2(_1235_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4267_ (.I(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4268_ (.A1(_1225_),
    .A2(_1230_),
    .B(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4269_ (.A1(_0988_),
    .A2(_0990_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4270_ (.A1(_1004_),
    .A2(_1238_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4271_ (.A1(_0908_),
    .A2(_0910_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4272_ (.I(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4273_ (.I(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4274_ (.A1(_1239_),
    .A2(_1004_),
    .A3(_1238_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4275_ (.A1(_1240_),
    .A2(_1243_),
    .A3(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4276_ (.I(_0940_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4277_ (.I(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4278_ (.A1(_1033_),
    .A2(_1049_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4279_ (.I(_1094_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4280_ (.A1(_3245_),
    .A2(_0896_),
    .A3(_0898_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4281_ (.I(_0574_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(_1250_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4283_ (.I(_0591_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4284_ (.A1(_1253_),
    .A2(_1093_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4285_ (.A1(_1249_),
    .A2(_1252_),
    .B(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4286_ (.A1(\mod.pc_2[6] ),
    .A2(_1205_),
    .B1(_0510_),
    .B2(_0523_),
    .C(_1047_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4287_ (.A1(_0551_),
    .A2(_1022_),
    .A3(_1026_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4288_ (.A1(_1033_),
    .A2(_1256_),
    .B(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4289_ (.A1(_1248_),
    .A2(_1255_),
    .B(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4290_ (.A1(_1062_),
    .A2(_1063_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4291_ (.A1(_0807_),
    .A2(_0650_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_0723_),
    .A2(_0666_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4293_ (.A1(_1260_),
    .A2(_1261_),
    .B(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4294_ (.A1(_0625_),
    .A2(_0680_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4295_ (.A1(_0578_),
    .A2(_0494_),
    .A3(_1069_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4296_ (.A1(_1265_),
    .A2(_1070_),
    .B1(_0460_),
    .B2(_0452_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4297_ (.A1(_1055_),
    .A2(_1061_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4298_ (.A1(_1264_),
    .A2(_1266_),
    .B(_1267_),
    .C(_1260_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4299_ (.A1(_0899_),
    .A2(_1251_),
    .B(_1075_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4300_ (.A1(_1033_),
    .A2(_1048_),
    .A3(_1094_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4301_ (.A1(_1263_),
    .A2(_1268_),
    .B(_1269_),
    .C(_1270_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4302_ (.A1(_1165_),
    .A2(_1166_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4303_ (.A1(_1180_),
    .A2(_1181_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4304_ (.A1(_1272_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4305_ (.A1(_1127_),
    .A2(_1150_),
    .A3(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4306_ (.A1(_1259_),
    .A2(_1271_),
    .B(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4307_ (.A1(_1161_),
    .A2(_1164_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4308_ (.A1(_0840_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4309_ (.A1(_0873_),
    .A2(_1124_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4310_ (.A1(_0859_),
    .A2(_1144_),
    .A3(_1146_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4311_ (.A1(_0874_),
    .A2(_1121_),
    .A3(_1123_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4312_ (.A1(_1279_),
    .A2(_1280_),
    .B(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4313_ (.A1(_1177_),
    .A2(_1179_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4314_ (.A1(_0826_),
    .A2(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4315_ (.A1(_1182_),
    .A2(_1278_),
    .B1(_1282_),
    .B2(_1274_),
    .C(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4316_ (.I(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4317_ (.A1(_1276_),
    .A2(_1286_),
    .B(_1223_),
    .C(_1203_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_1226_),
    .A2(_1202_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4319_ (.A1(_0731_),
    .A2(_0734_),
    .A3(_0737_),
    .A4(_0739_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4320_ (.A1(_0742_),
    .A2(_0744_),
    .A3(_0750_),
    .A4(_0753_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4321_ (.A1(\mod.pc_2[12] ),
    .A2(_1205_),
    .B1(_1289_),
    .B2(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4322_ (.A1(_1291_),
    .A2(_1220_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(_1203_),
    .A2(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4324_ (.A1(_1288_),
    .A2(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4325_ (.I(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4326_ (.A1(_1287_),
    .A2(_1295_),
    .B(_1236_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4327_ (.A1(_1003_),
    .A2(_1232_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4328_ (.A1(_1296_),
    .A2(_1297_),
    .B(_0992_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4329_ (.A1(_0991_),
    .A2(_1296_),
    .A3(_1297_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4330_ (.I(_0911_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4331_ (.I(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4332_ (.I(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4333_ (.A1(_1298_),
    .A2(_1299_),
    .B(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4334_ (.A1(_1298_),
    .A2(_1299_),
    .B(_3241_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4335_ (.I(_0808_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4336_ (.I(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4337_ (.I(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4338_ (.A1(_0683_),
    .A2(_0684_),
    .B(_0680_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4339_ (.A1(_0454_),
    .A2(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4340_ (.I(_1059_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4341_ (.A1(_0757_),
    .A2(_0861_),
    .A3(_0650_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4342_ (.A1(_0527_),
    .A2(_1310_),
    .B(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4343_ (.I(_0923_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4344_ (.I0(_1309_),
    .I1(_1312_),
    .S(_1313_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4345_ (.I(_0809_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4346_ (.I(_0801_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4347_ (.I(_1316_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4348_ (.A1(_0828_),
    .A2(_0861_),
    .B(_1253_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4349_ (.A1(_1074_),
    .A2(_0527_),
    .A3(_0573_),
    .B(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4350_ (.A1(_0757_),
    .A2(_0861_),
    .B(_0551_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4351_ (.A1(_0579_),
    .A2(_0525_),
    .A3(_0681_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4352_ (.A1(_1320_),
    .A2(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4353_ (.A1(_1317_),
    .A2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4354_ (.A1(_1317_),
    .A2(_1319_),
    .B(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4355_ (.A1(_1315_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4356_ (.A1(_1307_),
    .A2(_1314_),
    .B(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4357_ (.I(_0716_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4358_ (.I(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4359_ (.I(_0920_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_1328_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4361_ (.I(_0917_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4362_ (.I(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4363_ (.I(_0692_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4364_ (.A1(_1205_),
    .A2(_0799_),
    .A3(_3262_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4365_ (.A1(_1333_),
    .A2(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4366_ (.A1(_0878_),
    .A2(_1241_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4367_ (.I(_1250_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_1337_),
    .A2(_0724_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4369_ (.A1(_1336_),
    .A2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4370_ (.I(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4371_ (.I(_0621_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4372_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4373_ (.I(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4374_ (.I(_0625_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4375_ (.A1(_1344_),
    .A2(_0527_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4376_ (.A1(_1343_),
    .A2(_1345_),
    .B(_1336_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4377_ (.A1(_1328_),
    .A2(_1335_),
    .B(_1340_),
    .C(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(_1332_),
    .A2(_1347_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4379_ (.A1(_3229_),
    .A2(_3244_),
    .A3(_3247_),
    .A4(_0936_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4380_ (.I(_0621_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4381_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4383_ (.A1(_0926_),
    .A2(_0774_),
    .B(_0874_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4384_ (.A1(_0683_),
    .A2(_0684_),
    .A3(_0859_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4385_ (.A1(_1353_),
    .A2(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4386_ (.A1(_0813_),
    .A2(_0814_),
    .B(_0826_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4387_ (.I(_0460_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4388_ (.A1(_1357_),
    .A2(_0840_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4389_ (.A1(_1356_),
    .A2(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4390_ (.I0(_1355_),
    .I1(_1359_),
    .S(_0497_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4391_ (.A1(_1352_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4392_ (.A1(_0789_),
    .A2(_0813_),
    .A3(_0814_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4393_ (.A1(_0925_),
    .A2(_1334_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4394_ (.A1(_0529_),
    .A2(_1291_),
    .A3(_0553_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4395_ (.A1(_1226_),
    .A2(_1357_),
    .B(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4396_ (.A1(_0725_),
    .A2(_0920_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4397_ (.I(_1366_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4398_ (.A1(_1362_),
    .A2(_1363_),
    .B1(_1365_),
    .B2(_0627_),
    .C(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4399_ (.I(_0934_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4400_ (.A1(_0932_),
    .A2(_0936_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4401_ (.I(_1370_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4402_ (.A1(_0988_),
    .A2(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4403_ (.A1(_0990_),
    .A2(_1369_),
    .B(_1372_),
    .C(_1246_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4404_ (.A1(_0992_),
    .A2(_1349_),
    .B1(_1361_),
    .B2(_1368_),
    .C(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4405_ (.A1(_1326_),
    .A2(_1330_),
    .B(_1348_),
    .C(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4406_ (.A1(_1245_),
    .A2(_1247_),
    .A3(_1303_),
    .B1(_1304_),
    .B2(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4407_ (.I(_1376_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4408_ (.I(_0987_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4409_ (.A1(_0950_),
    .A2(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4410_ (.A1(_0992_),
    .A2(_1377_),
    .B(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4411_ (.A1(_0943_),
    .A2(_1377_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4412_ (.A1(_0942_),
    .A2(_0932_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4413_ (.I(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4414_ (.I(_1383_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4415_ (.I(_1384_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4416_ (.A1(_0943_),
    .A2(_1380_),
    .B(_1381_),
    .C(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4417_ (.A1(_0949_),
    .A2(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4418_ (.I(\mod.valid2 ),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4419_ (.I(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4420_ (.I(_3227_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4421_ (.I(_3229_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4422_ (.I(_0914_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4423_ (.A1(_1391_),
    .A2(_1380_),
    .B(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4424_ (.I(_1376_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4425_ (.A1(_0992_),
    .A2(_1394_),
    .B(_1391_),
    .C(_1379_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4426_ (.I(_1237_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4427_ (.I(_0945_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4428_ (.A1(_1396_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4429_ (.A1(_1237_),
    .A2(_1287_),
    .A3(_1295_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4430_ (.I(_0726_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_0667_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4432_ (.A1(_1401_),
    .A2(_1310_),
    .B(_0576_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4433_ (.A1(_0525_),
    .A2(_0461_),
    .B(_0592_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4434_ (.I0(_1402_),
    .I1(_1403_),
    .S(_1313_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4435_ (.A1(_0461_),
    .A2(_1054_),
    .B(_0682_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4436_ (.I(_0801_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4437_ (.I0(_1405_),
    .I1(_0462_),
    .S(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4438_ (.I0(_1404_),
    .I1(_1407_),
    .S(_1351_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4439_ (.A1(_0757_),
    .A2(_0774_),
    .B(_1291_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4440_ (.A1(_1409_),
    .A2(_0827_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4441_ (.A1(_0790_),
    .A2(_0775_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4442_ (.A1(_0627_),
    .A2(_1410_),
    .B1(_1411_),
    .B2(_1333_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4443_ (.A1(_0554_),
    .A2(_0860_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4444_ (.A1(_1357_),
    .A2(_0840_),
    .B(_0875_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4445_ (.I0(_1413_),
    .I1(_1414_),
    .S(_1313_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4446_ (.A1(_1351_),
    .A2(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4447_ (.A1(_1400_),
    .A2(_1412_),
    .A3(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4448_ (.A1(_1400_),
    .A2(_1408_),
    .B(_1417_),
    .C(_1329_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4449_ (.I(_0715_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4450_ (.I(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4451_ (.A1(_0924_),
    .A2(_0790_),
    .A3(_0800_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4452_ (.A1(_0923_),
    .A2(_1305_),
    .B(_0950_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4453_ (.A1(_1242_),
    .A2(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4454_ (.A1(_1420_),
    .A2(_1421_),
    .B(_1423_),
    .C(_1340_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4455_ (.A1(_1004_),
    .A2(_0934_),
    .B(_1246_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4456_ (.A1(_1235_),
    .A2(_1371_),
    .B1(_1424_),
    .B2(_1331_),
    .C(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4457_ (.A1(_1418_),
    .A2(_1426_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4458_ (.A1(_1296_),
    .A2(_3242_),
    .A3(_1399_),
    .B(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4459_ (.I(_1300_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4460_ (.A1(_1237_),
    .A2(_1225_),
    .A3(_1230_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4461_ (.A1(_1238_),
    .A2(_1429_),
    .A3(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4462_ (.I(_3250_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4463_ (.I(_1432_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4464_ (.A1(_1302_),
    .A2(_1296_),
    .A3(_1399_),
    .B(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4465_ (.A1(_1398_),
    .A2(_1428_),
    .B1(_1431_),
    .B2(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4466_ (.I(_1242_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4467_ (.I(_1097_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4468_ (.A1(_1253_),
    .A2(_1099_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4469_ (.A1(_1337_),
    .A2(_1251_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4470_ (.A1(_1253_),
    .A2(_1099_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4471_ (.A1(_1438_),
    .A2(_1439_),
    .B(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4472_ (.I(_1048_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4473_ (.A1(_1097_),
    .A2(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4474_ (.A1(_1437_),
    .A2(_1256_),
    .B1(_1441_),
    .B2(_1443_),
    .C(_1257_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4475_ (.A1(_1072_),
    .A2(_1063_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4476_ (.A1(_1341_),
    .A2(_1054_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4477_ (.A1(_0716_),
    .A2(_1310_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4478_ (.A1(_1445_),
    .A2(_1446_),
    .B(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4479_ (.A1(_0812_),
    .A2(_1069_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4480_ (.A1(_0688_),
    .A2(_0689_),
    .A3(_1069_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4481_ (.A1(_1068_),
    .A2(_1450_),
    .B(_0454_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4482_ (.A1(_1056_),
    .A2(_1061_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4483_ (.A1(_1449_),
    .A2(_1451_),
    .B(_1452_),
    .C(_1445_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4484_ (.I(_1269_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4485_ (.A1(_1097_),
    .A2(_1049_),
    .A3(_1249_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4486_ (.A1(_1448_),
    .A2(_1453_),
    .B(_1454_),
    .C(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4487_ (.A1(_1128_),
    .A2(_1151_),
    .A3(_1274_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4488_ (.A1(_1444_),
    .A2(_1456_),
    .B(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4489_ (.A1(_1228_),
    .A2(_1222_),
    .B1(_1458_),
    .B2(_1285_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4490_ (.A1(_1224_),
    .A2(_1276_),
    .A3(_1286_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4491_ (.A1(_1459_),
    .A2(_1460_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4492_ (.A1(_1436_),
    .A2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4493_ (.A1(_1184_),
    .A2(_1190_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4494_ (.A1(_1224_),
    .A2(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4495_ (.A1(_1302_),
    .A2(_1464_),
    .B(_1246_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4496_ (.A1(_3242_),
    .A2(_1461_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4497_ (.I(_0726_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(_0691_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4499_ (.A1(_1468_),
    .A2(_1305_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4500_ (.I0(_1403_),
    .I1(_1413_),
    .S(_0496_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4501_ (.A1(_0925_),
    .A2(_1410_),
    .B1(_1414_),
    .B2(_1469_),
    .C1(_1470_),
    .C2(_1315_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4502_ (.A1(_1467_),
    .A2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4503_ (.I(_0717_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4504_ (.A1(_0461_),
    .A2(_1054_),
    .B(_0682_),
    .C(_0923_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4505_ (.A1(_1401_),
    .A2(_1310_),
    .B(_0575_),
    .C(_0812_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4506_ (.A1(_1316_),
    .A2(_0927_),
    .B(_1350_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4507_ (.A1(_0811_),
    .A2(_1474_),
    .A3(_1475_),
    .B(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4508_ (.A1(_1473_),
    .A2(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4509_ (.A1(_1329_),
    .A2(_1472_),
    .A3(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4510_ (.A1(_0776_),
    .A2(_0803_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4511_ (.A1(_1351_),
    .A2(_1336_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4512_ (.A1(_1307_),
    .A2(_1480_),
    .B1(_1481_),
    .B2(_1337_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4513_ (.A1(_1473_),
    .A2(_1482_),
    .B(_1340_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4514_ (.I(_0937_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(_1484_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4516_ (.A1(_1228_),
    .A2(_1369_),
    .B(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4517_ (.A1(_1332_),
    .A2(_1483_),
    .B1(_1486_),
    .B2(_1222_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4518_ (.A1(_1224_),
    .A2(_1397_),
    .B(_1479_),
    .C(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4519_ (.A1(_1462_),
    .A2(_1465_),
    .B(_1466_),
    .C(_1488_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4520_ (.A1(_1148_),
    .A2(_1149_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4521_ (.A1(_1102_),
    .A2(_1105_),
    .A3(_1490_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4522_ (.I(_1490_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4523_ (.A1(_1102_),
    .A2(_1105_),
    .B(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4524_ (.A1(_1491_),
    .A2(_1493_),
    .B(_1242_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4525_ (.I(_0912_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4526_ (.A1(_1259_),
    .A2(_1271_),
    .B(_1151_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4527_ (.A1(_1492_),
    .A2(_1444_),
    .A3(_1456_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4528_ (.A1(_1495_),
    .A2(_1496_),
    .A3(_1497_),
    .B(_1432_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4529_ (.A1(_1496_),
    .A2(_1497_),
    .B(_1383_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4530_ (.A1(_1474_),
    .A2(_1475_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4531_ (.I(_1305_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4532_ (.I0(_1500_),
    .I1(_1470_),
    .S(_1501_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4533_ (.A1(_0924_),
    .A2(_0927_),
    .B(_0717_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4534_ (.A1(_1420_),
    .A2(_1502_),
    .B(_1503_),
    .C(_0920_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4535_ (.A1(_1327_),
    .A2(_0810_),
    .A3(_0877_),
    .B(_1339_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4536_ (.I(_1148_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4537_ (.A1(_1506_),
    .A2(_1349_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4538_ (.A1(_1506_),
    .A2(_0934_),
    .B(_1507_),
    .C(_1484_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4539_ (.A1(_0918_),
    .A2(_1505_),
    .B1(_1508_),
    .B2(_1149_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4540_ (.A1(_1504_),
    .A2(_1509_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4541_ (.A1(_1494_),
    .A2(_1498_),
    .B(_1499_),
    .C(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4542_ (.A1(_1448_),
    .A2(_1453_),
    .B(_1454_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4543_ (.A1(_1512_),
    .A2(_1439_),
    .B(_1438_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4544_ (.I(_1269_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4545_ (.A1(_1263_),
    .A2(_1268_),
    .B(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4546_ (.A1(_1249_),
    .A2(_1515_),
    .A3(_1252_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4547_ (.A1(_1513_),
    .A2(_1516_),
    .B(_1301_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_1073_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4549_ (.A1(_1518_),
    .A2(_1514_),
    .B(_1075_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4550_ (.A1(_1438_),
    .A2(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4551_ (.A1(_1438_),
    .A2(_1519_),
    .B(_1495_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4552_ (.A1(_1520_),
    .A2(_1521_),
    .B(_1432_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4553_ (.A1(_1383_),
    .A2(_1513_),
    .A3(_1516_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4554_ (.A1(_1344_),
    .A2(_1356_),
    .A3(_1364_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4555_ (.A1(_0529_),
    .A2(_0681_),
    .A3(_0839_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4556_ (.A1(_0593_),
    .A2(_1353_),
    .A3(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4557_ (.A1(_1524_),
    .A2(_1526_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4558_ (.A1(_1318_),
    .A2(_1321_),
    .B(_1406_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4559_ (.A1(_1320_),
    .A2(_1354_),
    .B(_1344_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4560_ (.A1(_0811_),
    .A2(_1528_),
    .A3(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4561_ (.A1(_1342_),
    .A2(_1527_),
    .B(_1530_),
    .C(_1419_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4562_ (.A1(_0691_),
    .A2(_1334_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4563_ (.A1(_0828_),
    .A2(_0553_),
    .B(_0773_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4564_ (.A1(_1362_),
    .A2(_1533_),
    .B(_0812_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4565_ (.A1(_1532_),
    .A2(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4566_ (.A1(_1501_),
    .A2(_1419_),
    .A3(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4567_ (.A1(_1401_),
    .A2(_0623_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(_0899_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4569_ (.A1(_1538_),
    .A2(_0724_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4570_ (.A1(_0989_),
    .A2(_1538_),
    .B1(_1422_),
    .B2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4571_ (.A1(_1241_),
    .A2(_1338_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4572_ (.A1(_0900_),
    .A2(_1537_),
    .B(_1540_),
    .C(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4573_ (.A1(_1531_),
    .A2(_1536_),
    .A3(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4574_ (.I0(_1312_),
    .I1(_1319_),
    .S(_0593_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4575_ (.A1(_1468_),
    .A2(_1501_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4576_ (.A1(_1306_),
    .A2(_1544_),
    .B1(_1545_),
    .B2(_1309_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4577_ (.A1(_1076_),
    .A2(_1099_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4578_ (.A1(_0930_),
    .A2(_0932_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4579_ (.I(_1548_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4580_ (.A1(_1547_),
    .A2(_0944_),
    .B(_0938_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4581_ (.A1(_1547_),
    .A2(_1549_),
    .B1(_1550_),
    .B2(_1098_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4582_ (.A1(_1367_),
    .A2(_1546_),
    .B(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4583_ (.A1(_1331_),
    .A2(_1543_),
    .B(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4584_ (.A1(_1517_),
    .A2(_1522_),
    .B(_1523_),
    .C(_1553_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4585_ (.A1(_1265_),
    .A2(_1070_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4586_ (.A1(_1555_),
    .A2(_0454_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4587_ (.A1(_1401_),
    .A2(_0912_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4588_ (.A1(_1556_),
    .A2(_1557_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4589_ (.A1(_1528_),
    .A2(_1529_),
    .B(_1342_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4590_ (.A1(_1308_),
    .A2(_1311_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4591_ (.I0(_0666_),
    .I1(_1251_),
    .S(_0667_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4592_ (.A1(_0692_),
    .A2(_1560_),
    .B1(_1561_),
    .B2(_0626_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4593_ (.A1(_1559_),
    .A2(_1562_),
    .B(_1327_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4594_ (.A1(_0989_),
    .A2(_1316_),
    .A3(_1341_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4595_ (.A1(_1357_),
    .A2(_1564_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4596_ (.I(_1541_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4597_ (.A1(_0901_),
    .A2(_1565_),
    .B(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4598_ (.A1(_1524_),
    .A2(_1526_),
    .B(_0623_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4599_ (.A1(_0809_),
    .A2(_1532_),
    .A3(_1534_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4600_ (.A1(_0726_),
    .A2(_1568_),
    .A3(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4601_ (.A1(_1563_),
    .A2(_1567_),
    .A3(_1570_),
    .B(_0918_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4602_ (.I(_1382_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4603_ (.A1(_1309_),
    .A2(_1333_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4604_ (.A1(_1068_),
    .A2(_0933_),
    .B(_0939_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4605_ (.A1(_1555_),
    .A2(_1349_),
    .B1(_1371_),
    .B2(_1450_),
    .C(_1574_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4606_ (.A1(_1366_),
    .A2(_1573_),
    .B(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4607_ (.A1(_1572_),
    .A2(_1556_),
    .B(_1576_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4608_ (.A1(_3250_),
    .A2(_1558_),
    .B1(_1571_),
    .B2(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4609_ (.A1(_0948_),
    .A2(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4610_ (.A1(_1449_),
    .A2(_1451_),
    .B(_1452_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4611_ (.A1(_1267_),
    .A2(_1264_),
    .A3(_1266_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4612_ (.A1(_1580_),
    .A2(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4613_ (.A1(_1071_),
    .A2(_1452_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_0912_),
    .A2(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4615_ (.A1(_1300_),
    .A2(_1582_),
    .B(_1584_),
    .C(_3250_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4616_ (.A1(_1572_),
    .A2(_1582_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4617_ (.A1(_1306_),
    .A2(_1407_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_1056_),
    .A2(_1549_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4619_ (.A1(_0938_),
    .A2(_1588_),
    .B(_1061_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4620_ (.A1(_1267_),
    .A2(_1349_),
    .B1(_0921_),
    .B2(_1587_),
    .C(_1589_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4621_ (.A1(_0827_),
    .A2(_0841_),
    .B(_0802_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4622_ (.A1(_0529_),
    .A2(_0773_),
    .A3(_0681_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4623_ (.A1(_1409_),
    .A2(_1592_),
    .B(_1344_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4624_ (.A1(_0691_),
    .A2(_0808_),
    .A3(_0790_),
    .A4(_0800_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4625_ (.A1(_1350_),
    .A2(_1591_),
    .A3(_1593_),
    .B(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4626_ (.A1(_1327_),
    .A2(_1595_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4627_ (.A1(_0593_),
    .A2(_0860_),
    .A3(_0875_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4628_ (.A1(_1313_),
    .A2(_0555_),
    .B(_1597_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4629_ (.A1(_0576_),
    .A2(_0592_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4630_ (.A1(_1469_),
    .A2(_1599_),
    .B1(_0668_),
    .B2(_0924_),
    .C(_0725_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4631_ (.A1(_1342_),
    .A2(_1598_),
    .B(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4632_ (.A1(_0901_),
    .A2(_1564_),
    .B(_1566_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4633_ (.A1(_1596_),
    .A2(_1601_),
    .A3(_1602_),
    .B(_0917_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4634_ (.A1(_1585_),
    .A2(_1586_),
    .A3(_1590_),
    .A4(_1603_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4635_ (.A1(_1300_),
    .A2(_0940_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4636_ (.A1(_1454_),
    .A2(_1448_),
    .A3(_1453_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4637_ (.A1(_1572_),
    .A2(_1605_),
    .B(_1606_),
    .C(_1515_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4638_ (.A1(_1316_),
    .A2(_0576_),
    .A3(_0592_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4639_ (.A1(_1468_),
    .A2(_0555_),
    .B(_1608_),
    .C(_0623_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4640_ (.A1(_0809_),
    .A2(_0842_),
    .A3(_0876_),
    .B(_0725_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4641_ (.A1(_0878_),
    .A2(_1341_),
    .A3(_0716_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4642_ (.A1(_0900_),
    .A2(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4643_ (.A1(_1501_),
    .A2(_1419_),
    .A3(_0776_),
    .A4(_0803_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4644_ (.A1(_1609_),
    .A2(_1610_),
    .B1(_1612_),
    .B2(_1566_),
    .C(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4645_ (.A1(_1518_),
    .A2(_1514_),
    .B(_1241_),
    .C(_0940_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4646_ (.A1(_1518_),
    .A2(_1269_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4647_ (.A1(_1074_),
    .A2(_1337_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4648_ (.A1(_1095_),
    .A2(_1370_),
    .B1(_1548_),
    .B2(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4649_ (.A1(_1514_),
    .A2(_0945_),
    .B1(_1366_),
    .B2(_1477_),
    .C(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4650_ (.A1(_0918_),
    .A2(_1614_),
    .B1(_1615_),
    .B2(_1616_),
    .C(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4651_ (.A1(_1607_),
    .A2(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4652_ (.A1(_1580_),
    .A2(_1261_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4653_ (.A1(_1445_),
    .A2(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4654_ (.A1(_1071_),
    .A2(_1267_),
    .B(_1056_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4655_ (.A1(_1260_),
    .A2(_1624_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4656_ (.A1(_1495_),
    .A2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4657_ (.A1(_1301_),
    .A2(_1623_),
    .B(_1626_),
    .C(_1432_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4658_ (.A1(_1320_),
    .A2(_1354_),
    .B(_1406_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4659_ (.A1(_1353_),
    .A2(_1525_),
    .B(_0496_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4660_ (.A1(_1628_),
    .A2(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4661_ (.A1(_1318_),
    .A2(_1321_),
    .A3(_0626_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4662_ (.A1(_0925_),
    .A2(_1561_),
    .B1(_1630_),
    .B2(_1306_),
    .C(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4663_ (.A1(_0989_),
    .A2(_1538_),
    .B(_1345_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4664_ (.A1(_1541_),
    .A2(_1612_),
    .A3(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4665_ (.A1(_1406_),
    .A2(_1362_),
    .A3(_1533_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4666_ (.A1(_0802_),
    .A2(_1356_),
    .A3(_1364_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4667_ (.A1(_1350_),
    .A2(_1334_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4668_ (.A1(_0811_),
    .A2(_1635_),
    .A3(_1636_),
    .B1(_1637_),
    .B2(_1468_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(_0717_),
    .A2(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4670_ (.A1(_1420_),
    .A2(_1632_),
    .B(_1634_),
    .C(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4671_ (.A1(_1315_),
    .A2(_1314_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4672_ (.A1(_1072_),
    .A2(_0944_),
    .B(_0938_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4673_ (.A1(_1072_),
    .A2(_1549_),
    .B1(_1642_),
    .B2(_1060_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4674_ (.A1(_1366_),
    .A2(_1641_),
    .B(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4675_ (.A1(_1572_),
    .A2(_1623_),
    .B1(_1640_),
    .B2(_1331_),
    .C(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4676_ (.A1(_1604_),
    .A2(_1621_),
    .A3(_1627_),
    .A4(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4677_ (.A1(_1511_),
    .A2(_1554_),
    .A3(_1579_),
    .A4(_1646_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4678_ (.I(_1280_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4679_ (.A1(_1259_),
    .A2(_1271_),
    .B(_1492_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4680_ (.A1(_1648_),
    .A2(_1649_),
    .B(_1128_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4681_ (.I(_1279_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4682_ (.A1(_1444_),
    .A2(_1456_),
    .B(_1151_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4683_ (.A1(_1651_),
    .A2(_1280_),
    .A3(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4684_ (.A1(_1650_),
    .A2(_1653_),
    .B(_1429_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4685_ (.A1(_1651_),
    .A2(_1506_),
    .A3(_1493_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4686_ (.A1(_1506_),
    .A2(_1493_),
    .B(_1651_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4687_ (.A1(_1243_),
    .A2(_1655_),
    .A3(_1656_),
    .B(_1433_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4688_ (.A1(_1383_),
    .A2(_1650_),
    .A3(_1653_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4689_ (.A1(_0942_),
    .A2(_0914_),
    .A3(_0915_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4690_ (.I(_1339_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4691_ (.A1(_1420_),
    .A2(_1568_),
    .A3(_1569_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4692_ (.A1(_1495_),
    .A2(_1338_),
    .A3(_1565_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4693_ (.A1(_1660_),
    .A2(_1661_),
    .A3(_1662_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4694_ (.A1(_1659_),
    .A2(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4695_ (.I(_1315_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4696_ (.I0(_1322_),
    .I1(_1355_),
    .S(_0497_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4697_ (.A1(_1307_),
    .A2(_1544_),
    .B(_0922_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4698_ (.A1(_1665_),
    .A2(_1666_),
    .B(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4699_ (.I(_0945_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4700_ (.I(_1549_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4701_ (.A1(_1126_),
    .A2(_1371_),
    .B1(_1670_),
    .B2(_1186_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4702_ (.A1(_1128_),
    .A2(_1669_),
    .B1(_1573_),
    .B2(_1330_),
    .C(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4703_ (.A1(_1664_),
    .A2(_1668_),
    .A3(_1672_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4704_ (.A1(_1654_),
    .A2(_1657_),
    .B(_1658_),
    .C(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4705_ (.A1(_0526_),
    .A2(_1103_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4706_ (.A1(_0526_),
    .A2(_1103_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4707_ (.A1(_1515_),
    .A2(_1252_),
    .B(_1249_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4708_ (.A1(_1675_),
    .A2(_1676_),
    .B1(_1440_),
    .B2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4709_ (.A1(_1442_),
    .A2(_1254_),
    .A3(_1513_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4710_ (.A1(_1678_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4711_ (.A1(_1098_),
    .A2(_1100_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4712_ (.A1(_1518_),
    .A2(_1096_),
    .B(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4713_ (.A1(_1442_),
    .A2(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4714_ (.A1(_1243_),
    .A2(_1683_),
    .B(_1433_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4715_ (.A1(_1436_),
    .A2(_1680_),
    .B(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4716_ (.A1(_1317_),
    .A2(_1409_),
    .A3(_1592_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4717_ (.A1(_0497_),
    .A2(_0827_),
    .A3(_0841_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4718_ (.A1(_1343_),
    .A2(_1686_),
    .A3(_1687_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4719_ (.A1(_1307_),
    .A2(_1598_),
    .B(_1688_),
    .C(_1328_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4720_ (.A1(_1467_),
    .A2(_1421_),
    .B1(_1540_),
    .B2(_1566_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4721_ (.A1(_1689_),
    .A2(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(_1675_),
    .A2(_1670_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4723_ (.A1(_1675_),
    .A2(_1669_),
    .B(_1484_),
    .C(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4724_ (.A1(_0526_),
    .A2(_1103_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4725_ (.A1(_0922_),
    .A2(_1408_),
    .B1(_1693_),
    .B2(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4726_ (.A1(_3242_),
    .A2(_1680_),
    .B1(_1691_),
    .B2(_1659_),
    .C(_1695_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4727_ (.A1(_1647_),
    .A2(_1674_),
    .A3(_1685_),
    .A4(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4728_ (.A1(_1435_),
    .A2(_1489_),
    .A3(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4729_ (.I(_1429_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4730_ (.I(_1437_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4731_ (.A1(_1700_),
    .A2(_1256_),
    .A3(_1678_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4732_ (.A1(_1256_),
    .A2(_1678_),
    .B(_1700_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4733_ (.A1(_1442_),
    .A2(_1682_),
    .B(_1675_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4734_ (.A1(_1437_),
    .A2(_1703_),
    .B(_1243_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4735_ (.A1(_1437_),
    .A2(_1703_),
    .B(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4736_ (.A1(_1699_),
    .A2(_1701_),
    .A3(_1702_),
    .B(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4737_ (.A1(_1701_),
    .A2(_1702_),
    .B(_1384_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4738_ (.A1(_1429_),
    .A2(_0901_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_1635_),
    .A2(_1636_),
    .B(_1343_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4740_ (.A1(_1352_),
    .A2(_1630_),
    .B(_1709_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4741_ (.A1(_1328_),
    .A2(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4742_ (.A1(_1346_),
    .A2(_1335_),
    .B(_1400_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4743_ (.A1(_1708_),
    .A2(_1711_),
    .A3(_1712_),
    .B(_1332_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4744_ (.A1(_1326_),
    .A2(_1367_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4745_ (.A1(_1030_),
    .A2(_1670_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4746_ (.I(_1031_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4747_ (.A1(_1030_),
    .A2(_1669_),
    .B(_1485_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4748_ (.A1(_1716_),
    .A2(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4749_ (.A1(_1713_),
    .A2(_1714_),
    .A3(_1715_),
    .A4(_1718_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4750_ (.A1(_1247_),
    .A2(_1706_),
    .B(_1707_),
    .C(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4751_ (.I(_1228_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4752_ (.A1(_1222_),
    .A2(_1463_),
    .B(_1721_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4753_ (.A1(_1722_),
    .A2(_1204_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4754_ (.A1(_1287_),
    .A2(_1293_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4755_ (.A1(_1204_),
    .A2(_1459_),
    .A3(_1292_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4756_ (.A1(_1724_),
    .A2(_1725_),
    .B(_1302_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4757_ (.A1(_1699_),
    .A2(_1723_),
    .B(_1726_),
    .C(_1247_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4758_ (.A1(_1724_),
    .A2(_1384_),
    .A3(_1725_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4759_ (.A1(_1538_),
    .A2(_1301_),
    .A3(_1537_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4760_ (.A1(_1665_),
    .A2(_1535_),
    .B1(_1729_),
    .B2(_1422_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_1473_),
    .A2(_1730_),
    .B(_1340_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4762_ (.A1(_1227_),
    .A2(_1485_),
    .B1(_1369_),
    .B2(_1229_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4763_ (.A1(_1333_),
    .A2(_1365_),
    .B1(_0627_),
    .B2(_1359_),
    .C1(_1666_),
    .C2(_1343_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4764_ (.A1(_0922_),
    .A2(_1733_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4765_ (.A1(_1204_),
    .A2(_1397_),
    .B1(_1546_),
    .B2(_1330_),
    .C(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4766_ (.A1(_1332_),
    .A2(_1731_),
    .B(_1732_),
    .C(_1735_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4767_ (.A1(_1728_),
    .A2(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4768_ (.I(_1281_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4769_ (.A1(_1280_),
    .A2(_1652_),
    .B(_1651_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4770_ (.A1(_1738_),
    .A2(_1739_),
    .B(_1167_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4771_ (.I(_1272_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4772_ (.A1(_1741_),
    .A2(_1281_),
    .A3(_1650_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4773_ (.A1(_1740_),
    .A2(_1742_),
    .B(_1699_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4774_ (.A1(_1102_),
    .A2(_1105_),
    .B(_1279_),
    .C(_1492_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4775_ (.A1(_1188_),
    .A2(_1744_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4776_ (.A1(_1741_),
    .A2(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4777_ (.A1(_1436_),
    .A2(_1746_),
    .B(_1433_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4778_ (.A1(_1384_),
    .A2(_1740_),
    .A3(_1742_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4779_ (.A1(_1165_),
    .A2(_1485_),
    .B1(_1369_),
    .B2(_1185_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4780_ (.A1(_1665_),
    .A2(_1415_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4781_ (.A1(_1352_),
    .A2(_1404_),
    .B(_1473_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4782_ (.A1(_1467_),
    .A2(_1587_),
    .B(_1329_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4783_ (.A1(_1750_),
    .A2(_1751_),
    .B(_1752_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4784_ (.A1(_1400_),
    .A2(_1595_),
    .B1(_1481_),
    .B2(_1317_),
    .C(_1660_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4785_ (.A1(_1167_),
    .A2(_1669_),
    .B1(_1754_),
    .B2(_1659_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4786_ (.A1(_1749_),
    .A2(_1753_),
    .A3(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4787_ (.A1(_1743_),
    .A2(_1747_),
    .B(_1748_),
    .C(_1756_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4788_ (.A1(_1720_),
    .A2(_1727_),
    .A3(_1737_),
    .A4(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4789_ (.A1(_1281_),
    .A2(_1650_),
    .B(_1741_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4790_ (.A1(_1278_),
    .A2(_1759_),
    .B(_1273_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4791_ (.A1(_1273_),
    .A2(_1278_),
    .A3(_1759_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4792_ (.A1(_1436_),
    .A2(_1760_),
    .A3(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4793_ (.A1(_1741_),
    .A2(_1745_),
    .B(_1166_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4794_ (.A1(_1273_),
    .A2(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4795_ (.A1(_1699_),
    .A2(_1764_),
    .B(_1247_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4796_ (.A1(_1760_),
    .A2(_1761_),
    .B(_3243_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4797_ (.A1(_1345_),
    .A2(_1481_),
    .B1(_1638_),
    .B2(_1467_),
    .C(_1660_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4798_ (.A1(_1352_),
    .A2(_1324_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4799_ (.A1(_1665_),
    .A2(_1360_),
    .B(_1367_),
    .C(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4800_ (.A1(_1181_),
    .A2(_1484_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4801_ (.A1(_1180_),
    .A2(_1670_),
    .B(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4802_ (.A1(_1182_),
    .A2(_1397_),
    .B1(_1641_),
    .B2(_1330_),
    .C(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4803_ (.A1(_1769_),
    .A2(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4804_ (.A1(_1659_),
    .A2(_1767_),
    .B(_1773_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4805_ (.A1(_1762_),
    .A2(_1765_),
    .B(_1766_),
    .C(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4806_ (.A1(_1394_),
    .A2(_1698_),
    .A3(_1758_),
    .A4(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4807_ (.A1(_1392_),
    .A2(_1395_),
    .A3(_1776_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4808_ (.A1(_1376_),
    .A2(_1698_),
    .A3(_1758_),
    .A4(_1775_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4809_ (.A1(_1390_),
    .A2(_1394_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4810_ (.A1(_1390_),
    .A2(_1778_),
    .B(_1779_),
    .C(_1392_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4811_ (.I(_0942_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4812_ (.A1(_1781_),
    .A2(_1394_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4813_ (.A1(_1390_),
    .A2(_1776_),
    .B(_1782_),
    .C(_0943_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _4814_ (.A1(_1390_),
    .A2(_1393_),
    .A3(_1777_),
    .B1(_1780_),
    .B2(_1783_),
    .B3(_1391_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4815_ (.A1(_0904_),
    .A2(_0905_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4816_ (.I(_1785_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4817_ (.A1(_0908_),
    .A2(_1784_),
    .B(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(_1787_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(_0902_),
    .A2(_1785_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4820_ (.I(_1789_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4821_ (.A1(_1790_),
    .A2(_1387_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_1191_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4823_ (.A1(_0903_),
    .A2(_0906_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4824_ (.A1(_1792_),
    .A2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4825_ (.A1(\mod.pc_2[0] ),
    .A2(_1078_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4826_ (.A1(_1794_),
    .A2(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _4827_ (.A1(_1389_),
    .A2(_1788_),
    .A3(_1791_),
    .A4(_1796_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4828_ (.A1(_1191_),
    .A2(_0907_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4829_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4830_ (.A1(net15),
    .A2(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4831_ (.A1(net14),
    .A2(_1798_),
    .B(_1800_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4832_ (.I(\mod.ldr_hzd[11] ),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4833_ (.A1(_1802_),
    .A2(_0429_),
    .B(_0632_),
    .C(_0846_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4834_ (.I(\mod.ldr_hzd[9] ),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4835_ (.I(_0633_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4836_ (.A1(_3275_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4837_ (.I(\mod.ldr_hzd[8] ),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4838_ (.I(_0637_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4839_ (.A1(_1808_),
    .A2(_0445_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4840_ (.I(\mod.ldr_hzd[10] ),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4841_ (.A1(_1804_),
    .A2(_1806_),
    .B1(_0661_),
    .B2(_1807_),
    .C1(_1809_),
    .C2(_1810_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4842_ (.I(\mod.ldr_hzd[0] ),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4843_ (.I(\mod.ldr_hzd[1] ),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4844_ (.I(\mod.ldr_hzd[2] ),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4845_ (.I(\mod.ldr_hzd[3] ),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4846_ (.I0(_1812_),
    .I1(_1813_),
    .I2(_1814_),
    .I3(_1815_),
    .S0(_1805_),
    .S1(_1808_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4847_ (.I(\mod.ldr_hzd[12] ),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4848_ (.I(\mod.ldr_hzd[13] ),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4849_ (.I(\mod.ldr_hzd[14] ),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4850_ (.I(\mod.ldr_hzd[15] ),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4851_ (.I0(_1817_),
    .I1(_1818_),
    .I2(_1819_),
    .I3(_1820_),
    .S0(_1805_),
    .S1(_1808_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4852_ (.I(\mod.ldr_hzd[6] ),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4853_ (.A1(_1822_),
    .A2(_1809_),
    .B(_0636_),
    .C(_0424_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4854_ (.I(\mod.ldr_hzd[5] ),
    .Z(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(\mod.ldr_hzd[4] ),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4856_ (.I(\mod.ldr_hzd[7] ),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4857_ (.A1(_1824_),
    .A2(_1806_),
    .B1(_0661_),
    .B2(_1825_),
    .C1(_0429_),
    .C2(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4858_ (.A1(_1823_),
    .A2(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4859_ (.A1(_0640_),
    .A2(_1816_),
    .B1(_1821_),
    .B2(_0848_),
    .C(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4860_ (.A1(_1803_),
    .A2(_1811_),
    .B(_1829_),
    .C(_3244_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4861_ (.A1(_1781_),
    .A2(_1191_),
    .A3(_0907_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4862_ (.I(_3213_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4863_ (.A1(_1817_),
    .A2(_1832_),
    .B(_0478_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4864_ (.I(_3160_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4865_ (.A1(_0480_),
    .A2(_3256_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4866_ (.A1(_1135_),
    .A2(_1136_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4867_ (.A1(_1820_),
    .A2(_1834_),
    .B1(_1835_),
    .B2(_1819_),
    .C1(_1836_),
    .C2(_1818_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4868_ (.A1(_1833_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4869_ (.A1(_1814_),
    .A2(_1835_),
    .B(_1015_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4870_ (.A1(_1815_),
    .A2(_1834_),
    .B1(_1836_),
    .B2(_1813_),
    .C1(_1812_),
    .C2(_1832_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4871_ (.A1(_1839_),
    .A2(_1840_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4872_ (.A1(_1824_),
    .A2(_1836_),
    .B(_0616_),
    .C(_0951_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4873_ (.A1(_1826_),
    .A2(_1834_),
    .B1(_1835_),
    .B2(_1822_),
    .C1(_1825_),
    .C2(_1832_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4874_ (.A1(_1807_),
    .A2(_1832_),
    .B(_1113_),
    .C(_0711_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _4875_ (.A1(_1802_),
    .A2(_1834_),
    .B1(_1835_),
    .B2(_1810_),
    .C1(_1836_),
    .C2(_1804_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4876_ (.A1(_1842_),
    .A2(_1843_),
    .B1(_1844_),
    .B2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4877_ (.A1(_1838_),
    .A2(_1841_),
    .A3(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4878_ (.I(\mod.instr_2[6] ),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4879_ (.I(_0490_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4880_ (.I(_3255_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4881_ (.A1(_1849_),
    .A2(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4882_ (.I(_1851_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4883_ (.A1(\mod.instr_2[4] ),
    .A2(_1850_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4885_ (.A1(\mod.ldr_hzd[3] ),
    .A2(_1852_),
    .B1(_1854_),
    .B2(\mod.ldr_hzd[1] ),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4886_ (.A1(\mod.instr_2[4] ),
    .A2(\mod.instr_2[3] ),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4887_ (.A1(_1849_),
    .A2(\mod.instr_2[3] ),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(_1857_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4889_ (.A1(\mod.ldr_hzd[0] ),
    .A2(_1856_),
    .B1(_1858_),
    .B2(\mod.ldr_hzd[2] ),
    .C(\mod.instr_2[5] ),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4890_ (.A1(_1855_),
    .A2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(\mod.instr_2[5] ),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4892_ (.I(_1856_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4893_ (.A1(\mod.ldr_hzd[4] ),
    .A2(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4894_ (.A1(\mod.ldr_hzd[6] ),
    .A2(_1858_),
    .B1(_1854_),
    .B2(\mod.ldr_hzd[5] ),
    .C1(_1851_),
    .C2(\mod.ldr_hzd[7] ),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4895_ (.A1(_1861_),
    .A2(_1863_),
    .A3(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4896_ (.A1(_1848_),
    .A2(_1860_),
    .A3(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4897_ (.A1(\mod.ldr_hzd[15] ),
    .A2(_1852_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4898_ (.A1(\mod.ldr_hzd[14] ),
    .A2(_1857_),
    .B1(_1853_),
    .B2(\mod.ldr_hzd[13] ),
    .C1(\mod.ldr_hzd[12] ),
    .C2(_1856_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4899_ (.A1(_1861_),
    .A2(_1867_),
    .A3(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4900_ (.A1(\mod.ldr_hzd[11] ),
    .A2(_1852_),
    .B1(_1854_),
    .B2(\mod.ldr_hzd[9] ),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4901_ (.A1(\mod.ldr_hzd[8] ),
    .A2(_1856_),
    .B1(_1858_),
    .B2(\mod.ldr_hzd[10] ),
    .C(\mod.instr_2[5] ),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4902_ (.A1(_1870_),
    .A2(_1871_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4903_ (.A1(\mod.instr_2[6] ),
    .A2(_1869_),
    .A3(_1872_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_1866_),
    .A2(_1873_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4905_ (.A1(_1831_),
    .A2(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4906_ (.A1(_1831_),
    .A2(_1847_),
    .B(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4907_ (.A1(_1802_),
    .A2(_1810_),
    .A3(_1804_),
    .A4(_1807_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4908_ (.A1(_1820_),
    .A2(_1819_),
    .A3(_1818_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4909_ (.A1(_1826_),
    .A2(_1822_),
    .A3(_1824_),
    .A4(_1825_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4910_ (.A1(_1815_),
    .A2(_1814_),
    .A3(_1813_),
    .A4(_1812_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4911_ (.A1(_1877_),
    .A2(_1878_),
    .A3(_1879_),
    .A4(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4912_ (.A1(_1830_),
    .A2(_1876_),
    .B1(_1881_),
    .B2(_1817_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4913_ (.A1(_1801_),
    .A2(_1882_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4914_ (.I(_1883_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4915_ (.I(_1788_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4916_ (.I(\mod.valid2 ),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4917_ (.A1(_1886_),
    .A2(_1883_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4918_ (.I(net13),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4919_ (.A1(_1885_),
    .A2(_1887_),
    .B(\mod.valid0 ),
    .C(_1888_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4920_ (.A1(_1884_),
    .A2(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4921_ (.I(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4922_ (.I(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4923_ (.I(\mod.pc[0] ),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4924_ (.A1(_1388_),
    .A2(_1787_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4925_ (.I(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_1895_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_1896_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4928_ (.A1(_1893_),
    .A2(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4929_ (.A1(_1884_),
    .A2(_1889_),
    .B(_1895_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4930_ (.I(_1899_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4931_ (.I(_1900_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4932_ (.A1(\mod.pc0[0] ),
    .A2(_1892_),
    .B1(_1898_),
    .B2(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4933_ (.A1(_1797_),
    .A2(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4934_ (.I(_3155_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4935_ (.A1(_3225_),
    .A2(_1387_),
    .B1(_1903_),
    .B2(_1904_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4936_ (.A1(_3224_),
    .A2(_1905_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4937_ (.A1(\mod.des.des_counter[0] ),
    .A2(_3150_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4938_ (.I(_1906_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4939_ (.I(_1907_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4940_ (.I(_3243_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4941_ (.A1(_1909_),
    .A2(_1578_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4942_ (.I(_1389_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4943_ (.I(_1787_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4944_ (.A1(_1911_),
    .A2(_1912_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4945_ (.I(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4946_ (.I(_1789_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_1789_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4948_ (.A1(_1206_),
    .A2(_3259_),
    .B(_1077_),
    .C(_3263_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4949_ (.A1(\mod.pc_2[1] ),
    .A2(_1046_),
    .A3(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4950_ (.A1(_1916_),
    .A2(_1918_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4951_ (.A1(_1915_),
    .A2(_1910_),
    .B(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4952_ (.I(\mod.pc0[1] ),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4953_ (.I(_1890_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4954_ (.I(_1900_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4955_ (.I(_1895_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4956_ (.I(_1924_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4957_ (.A1(\mod.pc[1] ),
    .A2(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4958_ (.A1(_1921_),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_1926_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4959_ (.A1(_1914_),
    .A2(_1920_),
    .B(_1927_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4960_ (.I(_3153_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4961_ (.A1(_0470_),
    .A2(_0488_),
    .B(_1929_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4962_ (.A1(_1908_),
    .A2(_1910_),
    .B1(_1928_),
    .B2(_0001_),
    .C(_1930_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4963_ (.A1(_0599_),
    .A2(_0613_),
    .B(_3223_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4964_ (.I(_1385_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4965_ (.A1(_1932_),
    .A2(_1604_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4966_ (.I(_1388_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(_1025_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4968_ (.A1(_3229_),
    .A2(_0954_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4969_ (.A1(_0954_),
    .A2(_0492_),
    .B(_1936_),
    .C(_0669_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4970_ (.A1(_1206_),
    .A2(_0492_),
    .B(_1045_),
    .C(_0669_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4971_ (.A1(_1917_),
    .A2(_1937_),
    .B(_1938_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4972_ (.A1(_1051_),
    .A2(_1935_),
    .A3(_1939_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4973_ (.A1(_1916_),
    .A2(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4974_ (.A1(_1915_),
    .A2(_1933_),
    .B(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4975_ (.A1(_1934_),
    .A2(_1912_),
    .A3(_1942_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4976_ (.I(\mod.pc[2] ),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4977_ (.A1(_1944_),
    .A2(_1897_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4978_ (.A1(\mod.pc0[2] ),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4979_ (.A1(_1943_),
    .A2(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4980_ (.A1(_3225_),
    .A2(_1933_),
    .B1(_1947_),
    .B2(_1904_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4981_ (.A1(_1931_),
    .A2(_1948_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4982_ (.A1(_0699_),
    .A2(_0710_),
    .B(_3223_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4983_ (.A1(_1627_),
    .A2(_1645_),
    .B(_1385_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4984_ (.I(_1145_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4985_ (.A1(_0651_),
    .A2(_1951_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4986_ (.A1(_1051_),
    .A2(_1935_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4987_ (.A1(_1051_),
    .A2(_1935_),
    .B1(_1917_),
    .B2(_1937_),
    .C(_1938_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4988_ (.A1(_1953_),
    .A2(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4989_ (.A1(_1952_),
    .A2(_1955_),
    .B(_1794_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4990_ (.A1(_1952_),
    .A2(_1955_),
    .B(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4991_ (.A1(_1915_),
    .A2(_1950_),
    .B(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4992_ (.A1(_1934_),
    .A2(_1788_),
    .A3(_1958_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4993_ (.I(_1890_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_1899_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4995_ (.I(\mod.pc[3] ),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4996_ (.I(_1924_),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4997_ (.A1(_1962_),
    .A2(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4998_ (.A1(\mod.pc0[3] ),
    .A2(_1960_),
    .B1(_1961_),
    .B2(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4999_ (.A1(_1959_),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5000_ (.A1(_3225_),
    .A2(_1950_),
    .B1(_1966_),
    .B2(_1904_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5001_ (.A1(_1949_),
    .A2(_1967_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5002_ (.A1(_1385_),
    .A2(_1621_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5003_ (.I(_3155_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5004_ (.I(_1794_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5005_ (.I(\mod.pc_2[4] ),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5006_ (.I(_1122_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5007_ (.A1(\mod.pc_2[3] ),
    .A2(_1951_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5008_ (.A1(\mod.pc_2[3] ),
    .A2(_1951_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5009_ (.A1(_1953_),
    .A2(_1973_),
    .A3(_1954_),
    .B(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5010_ (.A1(_1971_),
    .A2(_1972_),
    .A3(_1975_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5011_ (.A1(_1794_),
    .A2(_1968_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5012_ (.A1(_1970_),
    .A2(_1976_),
    .B(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5013_ (.A1(_1934_),
    .A2(_1912_),
    .A3(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5014_ (.I(\mod.pc[4] ),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5015_ (.A1(_1980_),
    .A2(_1897_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5016_ (.A1(\mod.pc0[4] ),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5017_ (.A1(_1979_),
    .A2(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5018_ (.A1(_1969_),
    .A2(_1983_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5019_ (.I(_3153_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5020_ (.A1(_0886_),
    .A2(_0895_),
    .B(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5021_ (.A1(_1908_),
    .A2(_1968_),
    .B(_1984_),
    .C(_1986_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5022_ (.I(_3154_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5023_ (.A1(_3243_),
    .A2(_1554_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5024_ (.A1(_1987_),
    .A2(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5025_ (.A1(_1082_),
    .A2(_1087_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(_1163_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5027_ (.A1(\mod.pc_2[4] ),
    .A2(_1972_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5028_ (.A1(_1971_),
    .A2(_1972_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5029_ (.A1(_1992_),
    .A2(_1975_),
    .B(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5030_ (.A1(\mod.pc_2[5] ),
    .A2(_1991_),
    .A3(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5031_ (.A1(_1916_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5032_ (.A1(_1915_),
    .A2(_1988_),
    .B(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5033_ (.A1(_1934_),
    .A2(_1912_),
    .A3(_1997_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5034_ (.I(\mod.pc[5] ),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5035_ (.A1(_1999_),
    .A2(_1963_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5036_ (.A1(\mod.pc0[5] ),
    .A2(_1960_),
    .B1(_1961_),
    .B2(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(_1998_),
    .A2(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5038_ (.A1(_3223_),
    .A2(_1990_),
    .B1(_2002_),
    .B2(_1904_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5039_ (.A1(_1989_),
    .A2(_2003_),
    .ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5040_ (.I(_1787_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5041_ (.I(_1916_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5042_ (.A1(_1685_),
    .A2(_1696_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5043_ (.A1(_1932_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5044_ (.I(\mod.pc_2[6] ),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5045_ (.I(_1178_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5046_ (.A1(\mod.pc_2[5] ),
    .A2(_1991_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5047_ (.A1(_2010_),
    .A2(_1994_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5048_ (.A1(\mod.pc_2[5] ),
    .A2(_1991_),
    .B(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5049_ (.A1(_2008_),
    .A2(_2009_),
    .A3(_2012_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5050_ (.A1(_1790_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5051_ (.A1(_2005_),
    .A2(_2007_),
    .B(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5052_ (.A1(_1911_),
    .A2(_2004_),
    .A3(_2015_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5053_ (.I(\mod.pc[6] ),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5054_ (.A1(_2017_),
    .A2(_1963_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5055_ (.A1(\mod.pc0[6] ),
    .A2(_1960_),
    .B1(_1961_),
    .B2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5056_ (.A1(_2016_),
    .A2(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5057_ (.A1(_1969_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5058_ (.A1(_1987_),
    .A2(_2007_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5059_ (.A1(_1037_),
    .A2(_1042_),
    .B(_1985_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5060_ (.A1(_2021_),
    .A2(_2022_),
    .A3(_2023_),
    .ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5061_ (.A1(_1909_),
    .A2(_1720_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5062_ (.I(_1208_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5063_ (.A1(\mod.pc_2[6] ),
    .A2(_2009_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5064_ (.A1(_2008_),
    .A2(_2009_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5065_ (.A1(_2026_),
    .A2(_2012_),
    .B(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5066_ (.A1(\mod.pc_2[7] ),
    .A2(_2025_),
    .A3(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_1790_),
    .A2(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5068_ (.A1(_2005_),
    .A2(_2024_),
    .B(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5069_ (.A1(_1911_),
    .A2(_2004_),
    .A3(_2031_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5070_ (.I(\mod.pc[7] ),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5071_ (.A1(_2033_),
    .A2(_1963_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5072_ (.A1(\mod.pc0[7] ),
    .A2(_1960_),
    .B1(_1961_),
    .B2(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5073_ (.A1(_2032_),
    .A2(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5074_ (.A1(_1969_),
    .A2(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5075_ (.A1(_1987_),
    .A2(_2024_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5076_ (.A1(_1008_),
    .A2(_1020_),
    .B(_1985_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5077_ (.A1(_2037_),
    .A2(_2038_),
    .A3(_2039_),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5078_ (.A1(_1909_),
    .A2(_1511_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5079_ (.I(_1896_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5080_ (.A1(_1135_),
    .A2(_0954_),
    .B(_0957_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5081_ (.A1(_0530_),
    .A2(_2025_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5082_ (.A1(_0530_),
    .A2(_2025_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5083_ (.A1(_2043_),
    .A2(_2028_),
    .B(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5084_ (.A1(_0843_),
    .A2(_2042_),
    .A3(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5085_ (.A1(_1970_),
    .A2(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5086_ (.A1(_1970_),
    .A2(_2040_),
    .B(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5087_ (.A1(_2041_),
    .A2(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5088_ (.I(\mod.pc[8] ),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5089_ (.A1(_2050_),
    .A2(_1896_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5090_ (.A1(\mod.pc0[8] ),
    .A2(_1892_),
    .B1(_1901_),
    .B2(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5091_ (.A1(_2049_),
    .A2(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5092_ (.A1(_1131_),
    .A2(_1142_),
    .B(_1929_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5093_ (.A1(_1908_),
    .A2(_2040_),
    .B1(_2053_),
    .B2(_0001_),
    .C(_2054_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5094_ (.A1(_1909_),
    .A2(_1674_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_1970_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5096_ (.A1(\mod.pc_2[8] ),
    .A2(_2042_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(\mod.pc_2[8] ),
    .A2(_2042_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5098_ (.A1(_2057_),
    .A2(_2045_),
    .B(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5099_ (.A1(\mod.pc_2[9] ),
    .A2(_1233_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5100_ (.A1(\mod.pc_2[9] ),
    .A2(_1233_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_2060_),
    .A2(_2061_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5102_ (.A1(_2059_),
    .A2(_2062_),
    .B(_1790_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5103_ (.A1(_2059_),
    .A2(_2062_),
    .B(_2063_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5104_ (.A1(_2056_),
    .A2(_2055_),
    .B(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5105_ (.I(\mod.pc[9] ),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5106_ (.A1(\mod.pc0[9] ),
    .A2(_1891_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5107_ (.A1(_2066_),
    .A2(_1891_),
    .B(_2067_),
    .C(_2041_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5108_ (.A1(_2041_),
    .A2(_2065_),
    .B(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5109_ (.A1(_1109_),
    .A2(_1120_),
    .B(_1929_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5110_ (.A1(_1908_),
    .A2(_2055_),
    .B1(_2069_),
    .B2(_0001_),
    .C(_2070_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5111_ (.A1(_0000_),
    .A2(\mod.des.des_counter[1] ),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5112_ (.I(_2071_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5113_ (.A1(_1156_),
    .A2(_1160_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5114_ (.A1(_1743_),
    .A2(_1747_),
    .B(_1756_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5115_ (.I(\mod.pc_2[10] ),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5116_ (.A1(_2075_),
    .A2(_0958_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5117_ (.I(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5118_ (.A1(_2059_),
    .A2(_2061_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5119_ (.A1(_2060_),
    .A2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5120_ (.A1(_2077_),
    .A2(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5121_ (.A1(_2060_),
    .A2(_2078_),
    .A3(_2076_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5122_ (.A1(_2005_),
    .A2(_2081_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5123_ (.A1(_2056_),
    .A2(_2074_),
    .B1(_2080_),
    .B2(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5124_ (.A1(_1914_),
    .A2(_2083_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5125_ (.I(\mod.pc[10] ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5126_ (.A1(_2085_),
    .A2(_1897_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5127_ (.A1(\mod.pc0[10] ),
    .A2(_1922_),
    .B1(_1923_),
    .B2(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5128_ (.A1(_2084_),
    .A2(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5129_ (.A1(_3225_),
    .A2(_2074_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5130_ (.A1(_2072_),
    .A2(_2073_),
    .B1(_2088_),
    .B2(_3156_),
    .C(_2089_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5131_ (.A1(_1932_),
    .A2(_1775_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5132_ (.A1(_2056_),
    .A2(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5133_ (.I(_2005_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5134_ (.A1(\mod.pc_2[10] ),
    .A2(_0958_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5135_ (.A1(_2093_),
    .A2(_2080_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5136_ (.I(\mod.pc_2[11] ),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5137_ (.A1(\mod.funct7[0] ),
    .A2(_1206_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5138_ (.A1(_0957_),
    .A2(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5139_ (.A1(_2095_),
    .A2(_2097_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5140_ (.A1(_2094_),
    .A2(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(_2092_),
    .A2(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5142_ (.A1(_1924_),
    .A2(_2091_),
    .A3(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5143_ (.I(\mod.pc[11] ),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5144_ (.A1(_2102_),
    .A2(_2041_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5145_ (.A1(\mod.pc0[11] ),
    .A2(_1892_),
    .B1(_1901_),
    .B2(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5146_ (.A1(_2101_),
    .A2(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5147_ (.A1(_1171_),
    .A2(_1176_),
    .B(_1929_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5148_ (.A1(_1907_),
    .A2(_2090_),
    .B1(_2105_),
    .B2(_3156_),
    .C(_2106_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5149_ (.I(_1932_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5150_ (.A1(_2107_),
    .A2(_1489_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(_1987_),
    .A2(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5152_ (.A1(\mod.pc_2[11] ),
    .A2(_2097_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5153_ (.A1(_2094_),
    .A2(_2098_),
    .B(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5154_ (.A1(\mod.pc_2[12] ),
    .A2(_1089_),
    .A3(_2111_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5155_ (.A1(_2092_),
    .A2(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5156_ (.A1(_2092_),
    .A2(_2108_),
    .B(_2113_),
    .C(_1924_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5157_ (.I(\mod.pc[12] ),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5158_ (.A1(_2115_),
    .A2(_1925_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5159_ (.A1(\mod.pc0[12] ),
    .A2(_1891_),
    .B1(_1900_),
    .B2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5160_ (.A1(_2114_),
    .A2(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5161_ (.A1(_1985_),
    .A2(_1218_),
    .B1(_2118_),
    .B2(_1969_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5162_ (.A1(_2109_),
    .A2(_2119_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5163_ (.A1(_1196_),
    .A2(_1199_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5164_ (.A1(_1727_),
    .A2(_1737_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5165_ (.A1(_2107_),
    .A2(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5166_ (.I(_0727_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5167_ (.A1(_2123_),
    .A2(_1089_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5168_ (.A1(_2123_),
    .A2(_1089_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5169_ (.A1(_2124_),
    .A2(_2111_),
    .B(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5170_ (.A1(\mod.pc_2[13] ),
    .A2(_0955_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5171_ (.A1(_2126_),
    .A2(_2127_),
    .B(_2056_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5172_ (.A1(_2126_),
    .A2(_2127_),
    .B(_2128_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5173_ (.A1(_2092_),
    .A2(_2122_),
    .B(_2129_),
    .C(_1896_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5174_ (.I(\mod.pc[13] ),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5175_ (.A1(_2131_),
    .A2(_1925_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5176_ (.A1(\mod.pc0[13] ),
    .A2(_1892_),
    .B1(_1901_),
    .B2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5177_ (.A1(_2130_),
    .A2(_2133_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5178_ (.A1(_3154_),
    .A2(_2122_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5179_ (.A1(_2072_),
    .A2(_2120_),
    .B1(_2134_),
    .B2(_3156_),
    .C(_2135_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5180_ (.I(_2107_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5181_ (.A1(_1907_),
    .A2(_2136_),
    .A3(_1435_),
    .B1(_1001_),
    .B2(_2072_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5182_ (.A1(_1907_),
    .A2(_2136_),
    .A3(_1377_),
    .B1(_0984_),
    .B2(_2072_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5183_ (.A1(_1792_),
    .A2(_0907_),
    .A3(_1887_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5184_ (.I(_2137_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5185_ (.A1(_1781_),
    .A2(net31),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5186_ (.I(_2138_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5187_ (.I(net11),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5188_ (.I(_2139_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5189_ (.I(_2140_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5190_ (.I(_1861_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5191_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .A3(net15),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5192_ (.I(_2142_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5193_ (.I(_2142_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5194_ (.A1(\mod.rd_3[2] ),
    .A2(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5195_ (.A1(_2141_),
    .A2(_2143_),
    .B(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5196_ (.I(_1848_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5197_ (.A1(\mod.rd_3[3] ),
    .A2(_2144_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5198_ (.A1(_2147_),
    .A2(_2143_),
    .B(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5199_ (.A1(_2146_),
    .A2(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5200_ (.A1(net12),
    .A2(_1883_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5201_ (.A1(_1886_),
    .A2(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(net12),
    .A2(_2142_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5203_ (.A1(_3244_),
    .A2(_2152_),
    .B(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5204_ (.I(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5205_ (.A1(\mod.rd_3[1] ),
    .A2(_2144_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5206_ (.A1(_1849_),
    .A2(_2143_),
    .B(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5207_ (.A1(\mod.rd_3[0] ),
    .A2(_2144_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5208_ (.A1(_1850_),
    .A2(_2143_),
    .B(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5209_ (.I(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5210_ (.A1(_2155_),
    .A2(_2157_),
    .A3(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5211_ (.A1(_2150_),
    .A2(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5212_ (.I(_2162_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5213_ (.I(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5214_ (.I(_2142_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5215_ (.I(_2165_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5216_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5217_ (.I(_1786_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5218_ (.I(_1786_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5219_ (.A1(_2169_),
    .A2(_1387_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5220_ (.A1(\mod.ins_ldr_3 ),
    .A2(\mod.valid_out3 ),
    .A3(net15),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5221_ (.A1(_1792_),
    .A2(_3257_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(_2171_),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5223_ (.I(_2173_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5224_ (.A1(_3263_),
    .A2(_2168_),
    .B(_2170_),
    .C(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5225_ (.A1(\mod.des.des_dout[21] ),
    .A2(_2167_),
    .B(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5226_ (.I(_2176_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5227_ (.I(_2162_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5228_ (.I(_2178_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5229_ (.A1(\mod.registers.r1[0] ),
    .A2(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5230_ (.A1(_2164_),
    .A2(_2177_),
    .B(_2180_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5231_ (.I(_1793_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5232_ (.I(_1793_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5233_ (.A1(\mod.pc_2[1] ),
    .A2(_2182_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5234_ (.A1(_2181_),
    .A2(_1910_),
    .B(_2174_),
    .C(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5235_ (.A1(\mod.des.des_dout[22] ),
    .A2(_2167_),
    .B(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5236_ (.I(_2185_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(\mod.registers.r1[1] ),
    .A2(_2179_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5238_ (.A1(_2164_),
    .A2(_2186_),
    .B(_2187_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5239_ (.I(_2165_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5240_ (.I(_2182_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5241_ (.A1(_2136_),
    .A2(_1604_),
    .B(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5242_ (.I(_2169_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5243_ (.A1(_0628_),
    .A2(_2191_),
    .B(_2174_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5244_ (.A1(\mod.des.des_dout[23] ),
    .A2(_2188_),
    .B1(_2190_),
    .B2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5245_ (.I(_2193_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5246_ (.A1(\mod.registers.r1[2] ),
    .A2(_2179_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5247_ (.A1(_2164_),
    .A2(_2194_),
    .B(_2195_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5248_ (.A1(_2169_),
    .A2(_1950_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5249_ (.A1(_0651_),
    .A2(_2168_),
    .B(_2173_),
    .C(_2196_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5250_ (.A1(\mod.des.des_dout[24] ),
    .A2(_2167_),
    .B(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_2198_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(\mod.registers.r1[3] ),
    .A2(_2179_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5253_ (.A1(_2164_),
    .A2(_2199_),
    .B(_2200_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5254_ (.I(_2163_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5255_ (.A1(_1971_),
    .A2(_2182_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5256_ (.A1(_2181_),
    .A2(_1968_),
    .B(_2173_),
    .C(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5257_ (.A1(\mod.des.des_dout[25] ),
    .A2(_2167_),
    .B(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5258_ (.I(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5259_ (.I(_2178_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5260_ (.A1(\mod.registers.r1[4] ),
    .A2(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5261_ (.A1(_2201_),
    .A2(_2205_),
    .B(_2207_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5262_ (.I(_2172_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5263_ (.I(_2208_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5264_ (.I(_1793_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5265_ (.A1(_2210_),
    .A2(_1988_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5266_ (.A1(_0580_),
    .A2(_2189_),
    .B(_2209_),
    .C(_2211_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5267_ (.I(_2165_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5268_ (.I(_2172_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5269_ (.A1(_1078_),
    .A2(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5270_ (.A1(_2213_),
    .A2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5271_ (.A1(\mod.des.des_dout[26] ),
    .A2(_2188_),
    .B1(_2212_),
    .B2(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5272_ (.I(_2217_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5273_ (.A1(\mod.registers.r1[5] ),
    .A2(_2206_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5274_ (.A1(_2201_),
    .A2(_2218_),
    .B(_2219_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5275_ (.I(_2171_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5276_ (.I(_1786_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5277_ (.A1(_2221_),
    .A2(_2007_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5278_ (.A1(_2008_),
    .A2(_2210_),
    .B(_2208_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5279_ (.A1(_0902_),
    .A2(_0561_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5280_ (.A1(_1046_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5281_ (.I(_2171_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5282_ (.A1(_2222_),
    .A2(_2223_),
    .B(_2225_),
    .C(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5283_ (.A1(\mod.des.des_dout[27] ),
    .A2(_2220_),
    .B(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5284_ (.I(_2228_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5285_ (.A1(\mod.registers.r1[6] ),
    .A2(_2206_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5286_ (.A1(_2201_),
    .A2(_2229_),
    .B(_2230_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5287_ (.A1(_2181_),
    .A2(_2024_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5288_ (.A1(\mod.pc_2[7] ),
    .A2(_2221_),
    .B(_2224_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5289_ (.A1(_1935_),
    .A2(_2208_),
    .B(_2226_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5290_ (.A1(_2231_),
    .A2(_2232_),
    .B(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5291_ (.A1(\mod.des.des_dout[28] ),
    .A2(_2188_),
    .B(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5292_ (.I(_2235_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5293_ (.A1(\mod.registers.r1[7] ),
    .A2(_2206_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5294_ (.A1(_2201_),
    .A2(_2236_),
    .B(_2237_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5295_ (.I(_2163_),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(\mod.pc_2[8] ),
    .A2(_2221_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5297_ (.A1(_2191_),
    .A2(_2040_),
    .B(_2209_),
    .C(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5298_ (.I(_2208_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5299_ (.A1(_1951_),
    .A2(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5300_ (.A1(_2213_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5301_ (.A1(\mod.des.des_dout[29] ),
    .A2(_2188_),
    .B1(_2240_),
    .B2(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5302_ (.I(_2244_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5303_ (.I(_2178_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5304_ (.A1(\mod.registers.r1[8] ),
    .A2(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5305_ (.A1(_2238_),
    .A2(_2245_),
    .B(_2247_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5306_ (.I(_2165_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5307_ (.A1(\mod.pc_2[9] ),
    .A2(_2221_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5308_ (.A1(_2191_),
    .A2(_2055_),
    .B(_2209_),
    .C(_2249_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5309_ (.A1(_1972_),
    .A2(_2241_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5310_ (.A1(_2213_),
    .A2(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5311_ (.A1(\mod.des.des_dout[30] ),
    .A2(_2248_),
    .B1(_2250_),
    .B2(_2252_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_2253_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5313_ (.A1(\mod.registers.r1[9] ),
    .A2(_2246_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5314_ (.A1(_2238_),
    .A2(_2254_),
    .B(_2255_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5315_ (.A1(_2210_),
    .A2(_2074_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5316_ (.A1(_2075_),
    .A2(_2189_),
    .B(_2209_),
    .C(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(_1991_),
    .A2(_2226_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5318_ (.A1(_2174_),
    .A2(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5319_ (.A1(\mod.des.des_dout[31] ),
    .A2(_2248_),
    .B1(_2257_),
    .B2(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5320_ (.I(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5321_ (.A1(\mod.registers.r1[10] ),
    .A2(_2246_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5322_ (.A1(_2238_),
    .A2(_2261_),
    .B(_2262_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5323_ (.A1(\mod.pc_2[11] ),
    .A2(_2169_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5324_ (.A1(_2191_),
    .A2(_2090_),
    .B(_2214_),
    .C(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5325_ (.A1(_2009_),
    .A2(_2241_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5326_ (.A1(_2166_),
    .A2(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5327_ (.A1(\mod.des.des_dout[32] ),
    .A2(_2248_),
    .B1(_2264_),
    .B2(_2266_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(_2267_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5329_ (.A1(\mod.registers.r1[11] ),
    .A2(_2246_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5330_ (.A1(_2238_),
    .A2(_2268_),
    .B(_2269_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5331_ (.I(_2163_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5332_ (.A1(_2210_),
    .A2(_2108_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5333_ (.A1(_2123_),
    .A2(_2189_),
    .B(_2214_),
    .C(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5334_ (.I(_2224_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5335_ (.A1(_2025_),
    .A2(_2273_),
    .B(_2166_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5336_ (.A1(\mod.des.des_dout[33] ),
    .A2(_2248_),
    .B1(_2272_),
    .B2(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5337_ (.I(_2275_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5338_ (.I(_2178_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5339_ (.A1(\mod.registers.r1[12] ),
    .A2(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5340_ (.A1(_2270_),
    .A2(_2276_),
    .B(_2278_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5341_ (.A1(_2182_),
    .A2(_2122_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5342_ (.A1(_0758_),
    .A2(_2181_),
    .B(_2214_),
    .C(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5343_ (.A1(_2042_),
    .A2(_2241_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5344_ (.A1(_2166_),
    .A2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5345_ (.A1(\mod.des.des_dout[34] ),
    .A2(_2213_),
    .B1(_2280_),
    .B2(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5346_ (.I(_2283_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(\mod.registers.r1[13] ),
    .A2(_2277_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5348_ (.A1(_2270_),
    .A2(_2284_),
    .B(_2285_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5349_ (.A1(_2168_),
    .A2(_2136_),
    .A3(_1435_),
    .A4(_2273_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5350_ (.A1(_1233_),
    .A2(_2273_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(_2220_),
    .A2(_2287_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5352_ (.A1(\mod.des.des_dout[35] ),
    .A2(_2220_),
    .B1(_2286_),
    .B2(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_2289_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5354_ (.A1(\mod.registers.r1[14] ),
    .A2(_2277_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5355_ (.A1(_2270_),
    .A2(_2290_),
    .B(_2291_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5356_ (.A1(_2168_),
    .A2(_2107_),
    .A3(_1377_),
    .A4(_2273_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5357_ (.A1(_0958_),
    .A2(_2224_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5358_ (.A1(_2226_),
    .A2(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5359_ (.A1(\mod.des.des_dout[36] ),
    .A2(_2220_),
    .B1(_2292_),
    .B2(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5360_ (.I(_2295_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(\mod.registers.r1[15] ),
    .A2(_2277_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5362_ (.A1(_2270_),
    .A2(_2296_),
    .B(_2297_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5363_ (.A1(_2154_),
    .A2(_2157_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5364_ (.A1(_2159_),
    .A2(_2298_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(_2150_),
    .A2(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5366_ (.I(_2300_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5367_ (.I(_2301_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5368_ (.I(_2300_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5369_ (.I(_2303_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5370_ (.A1(\mod.registers.r2[0] ),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5371_ (.A1(_2177_),
    .A2(_2302_),
    .B(_2305_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5372_ (.A1(\mod.registers.r2[1] ),
    .A2(_2304_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5373_ (.A1(_2186_),
    .A2(_2302_),
    .B(_2306_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5374_ (.A1(\mod.registers.r2[2] ),
    .A2(_2304_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5375_ (.A1(_2194_),
    .A2(_2302_),
    .B(_2307_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5376_ (.A1(\mod.registers.r2[3] ),
    .A2(_2304_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5377_ (.A1(_2199_),
    .A2(_2302_),
    .B(_2308_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5378_ (.I(_2301_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5379_ (.I(_2303_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5380_ (.A1(\mod.registers.r2[4] ),
    .A2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5381_ (.A1(_2205_),
    .A2(_2309_),
    .B(_2311_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5382_ (.A1(\mod.registers.r2[5] ),
    .A2(_2310_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5383_ (.A1(_2218_),
    .A2(_2309_),
    .B(_2312_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5384_ (.A1(\mod.registers.r2[6] ),
    .A2(_2310_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5385_ (.A1(_2229_),
    .A2(_2309_),
    .B(_2313_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5386_ (.A1(\mod.registers.r2[7] ),
    .A2(_2310_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5387_ (.A1(_2236_),
    .A2(_2309_),
    .B(_2314_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5388_ (.I(_2301_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5389_ (.I(_2303_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5390_ (.A1(\mod.registers.r2[8] ),
    .A2(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5391_ (.A1(_2245_),
    .A2(_2315_),
    .B(_2317_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(\mod.registers.r2[9] ),
    .A2(_2316_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5393_ (.A1(_2254_),
    .A2(_2315_),
    .B(_2318_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5394_ (.A1(\mod.registers.r2[10] ),
    .A2(_2316_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5395_ (.A1(_2261_),
    .A2(_2315_),
    .B(_2319_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5396_ (.A1(\mod.registers.r2[11] ),
    .A2(_2316_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5397_ (.A1(_2268_),
    .A2(_2315_),
    .B(_2320_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5398_ (.I(_2301_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5399_ (.I(_2303_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5400_ (.A1(\mod.registers.r2[12] ),
    .A2(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5401_ (.A1(_2276_),
    .A2(_2321_),
    .B(_2323_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5402_ (.A1(\mod.registers.r2[13] ),
    .A2(_2322_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5403_ (.A1(_2284_),
    .A2(_2321_),
    .B(_2324_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(\mod.registers.r2[14] ),
    .A2(_2322_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5405_ (.A1(_2290_),
    .A2(_2321_),
    .B(_2325_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5406_ (.A1(\mod.registers.r2[15] ),
    .A2(_2322_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5407_ (.A1(_2296_),
    .A2(_2321_),
    .B(_2326_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5408_ (.A1(_2160_),
    .A2(_2298_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5409_ (.A1(_2150_),
    .A2(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5410_ (.I(_2328_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_2329_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5412_ (.I(_2328_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5413_ (.I(_2331_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5414_ (.A1(\mod.registers.r3[0] ),
    .A2(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5415_ (.A1(_2177_),
    .A2(_2330_),
    .B(_2333_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5416_ (.A1(\mod.registers.r3[1] ),
    .A2(_2332_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5417_ (.A1(_2186_),
    .A2(_2330_),
    .B(_2334_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5418_ (.A1(\mod.registers.r3[2] ),
    .A2(_2332_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5419_ (.A1(_2194_),
    .A2(_2330_),
    .B(_2335_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5420_ (.A1(\mod.registers.r3[3] ),
    .A2(_2332_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5421_ (.A1(_2199_),
    .A2(_2330_),
    .B(_2336_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5422_ (.I(_2329_),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5423_ (.I(_2331_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5424_ (.A1(\mod.registers.r3[4] ),
    .A2(_2338_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5425_ (.A1(_2205_),
    .A2(_2337_),
    .B(_2339_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5426_ (.A1(\mod.registers.r3[5] ),
    .A2(_2338_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5427_ (.A1(_2218_),
    .A2(_2337_),
    .B(_2340_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5428_ (.A1(\mod.registers.r3[6] ),
    .A2(_2338_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5429_ (.A1(_2229_),
    .A2(_2337_),
    .B(_2341_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5430_ (.A1(\mod.registers.r3[7] ),
    .A2(_2338_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5431_ (.A1(_2236_),
    .A2(_2337_),
    .B(_2342_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5432_ (.I(_2329_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5433_ (.I(_2331_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5434_ (.A1(\mod.registers.r3[8] ),
    .A2(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5435_ (.A1(_2245_),
    .A2(_2343_),
    .B(_2345_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5436_ (.A1(\mod.registers.r3[9] ),
    .A2(_2344_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5437_ (.A1(_2254_),
    .A2(_2343_),
    .B(_2346_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5438_ (.A1(\mod.registers.r3[10] ),
    .A2(_2344_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5439_ (.A1(_2261_),
    .A2(_2343_),
    .B(_2347_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5440_ (.A1(\mod.registers.r3[11] ),
    .A2(_2344_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5441_ (.A1(_2268_),
    .A2(_2343_),
    .B(_2348_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5442_ (.I(_2329_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5443_ (.I(_2331_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5444_ (.A1(\mod.registers.r3[12] ),
    .A2(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5445_ (.A1(_2276_),
    .A2(_2349_),
    .B(_2351_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5446_ (.A1(\mod.registers.r3[13] ),
    .A2(_2350_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5447_ (.A1(_2284_),
    .A2(_2349_),
    .B(_2352_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5448_ (.A1(\mod.registers.r3[14] ),
    .A2(_2350_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5449_ (.A1(_2290_),
    .A2(_2349_),
    .B(_2353_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5450_ (.A1(\mod.registers.r3[15] ),
    .A2(_2350_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5451_ (.A1(_2296_),
    .A2(_2349_),
    .B(_2354_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5452_ (.I(_2146_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5453_ (.A1(_2355_),
    .A2(_2149_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5454_ (.A1(_2155_),
    .A2(_2157_),
    .A3(_2159_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5455_ (.A1(_2356_),
    .A2(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5456_ (.I(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5457_ (.I(_2359_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5458_ (.I(_2358_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5460_ (.A1(\mod.registers.r4[0] ),
    .A2(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5461_ (.A1(_2177_),
    .A2(_2360_),
    .B(_2363_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5462_ (.A1(\mod.registers.r4[1] ),
    .A2(_2362_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5463_ (.A1(_2186_),
    .A2(_2360_),
    .B(_2364_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5464_ (.A1(\mod.registers.r4[2] ),
    .A2(_2362_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5465_ (.A1(_2194_),
    .A2(_2360_),
    .B(_2365_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5466_ (.A1(\mod.registers.r4[3] ),
    .A2(_2362_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5467_ (.A1(_2199_),
    .A2(_2360_),
    .B(_2366_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5468_ (.I(_2359_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_2361_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5470_ (.A1(\mod.registers.r4[4] ),
    .A2(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5471_ (.A1(_2205_),
    .A2(_2367_),
    .B(_2369_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5472_ (.A1(\mod.registers.r4[5] ),
    .A2(_2368_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5473_ (.A1(_2218_),
    .A2(_2367_),
    .B(_2370_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5474_ (.A1(\mod.registers.r4[6] ),
    .A2(_2368_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5475_ (.A1(_2229_),
    .A2(_2367_),
    .B(_2371_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5476_ (.A1(\mod.registers.r4[7] ),
    .A2(_2368_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5477_ (.A1(_2236_),
    .A2(_2367_),
    .B(_2372_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5478_ (.I(_2359_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5479_ (.I(_2361_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5480_ (.A1(\mod.registers.r4[8] ),
    .A2(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5481_ (.A1(_2245_),
    .A2(_2373_),
    .B(_2375_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5482_ (.A1(\mod.registers.r4[9] ),
    .A2(_2374_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5483_ (.A1(_2254_),
    .A2(_2373_),
    .B(_2376_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5484_ (.A1(\mod.registers.r4[10] ),
    .A2(_2374_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5485_ (.A1(_2261_),
    .A2(_2373_),
    .B(_2377_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5486_ (.A1(\mod.registers.r4[11] ),
    .A2(_2374_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5487_ (.A1(_2268_),
    .A2(_2373_),
    .B(_2378_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5488_ (.I(_2359_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5489_ (.I(_2361_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5490_ (.A1(\mod.registers.r4[12] ),
    .A2(_2380_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5491_ (.A1(_2276_),
    .A2(_2379_),
    .B(_2381_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5492_ (.A1(\mod.registers.r4[13] ),
    .A2(_2380_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5493_ (.A1(_2284_),
    .A2(_2379_),
    .B(_2382_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5494_ (.A1(\mod.registers.r4[14] ),
    .A2(_2380_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5495_ (.A1(_2290_),
    .A2(_2379_),
    .B(_2383_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5496_ (.A1(\mod.registers.r4[15] ),
    .A2(_2380_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5497_ (.A1(_2296_),
    .A2(_2379_),
    .B(_2384_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5498_ (.I(_2176_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5499_ (.I(_2385_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5500_ (.A1(_2161_),
    .A2(_2356_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5501_ (.I(_2387_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5502_ (.I(_2388_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5503_ (.I(_2387_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5504_ (.I(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5505_ (.A1(\mod.registers.r5[0] ),
    .A2(_2391_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5506_ (.A1(_2386_),
    .A2(_2389_),
    .B(_2392_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5507_ (.I(_2185_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5508_ (.I(_2393_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5509_ (.A1(\mod.registers.r5[1] ),
    .A2(_2391_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5510_ (.A1(_2394_),
    .A2(_2389_),
    .B(_2395_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5511_ (.I(_2193_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5512_ (.I(_2396_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5513_ (.A1(\mod.registers.r5[2] ),
    .A2(_2391_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5514_ (.A1(_2397_),
    .A2(_2389_),
    .B(_2398_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5515_ (.I(_2198_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5516_ (.I(_2399_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5517_ (.A1(\mod.registers.r5[3] ),
    .A2(_2391_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5518_ (.A1(_2400_),
    .A2(_2389_),
    .B(_2401_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5519_ (.I(_2204_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5520_ (.I(_2402_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5521_ (.I(_2388_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5522_ (.I(_2390_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5523_ (.A1(\mod.registers.r5[4] ),
    .A2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5524_ (.A1(_2403_),
    .A2(_2404_),
    .B(_2406_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5525_ (.I(_2217_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5526_ (.I(_2407_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5527_ (.A1(\mod.registers.r5[5] ),
    .A2(_2405_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5528_ (.A1(_2408_),
    .A2(_2404_),
    .B(_2409_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5529_ (.I(_2228_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5530_ (.I(_2410_),
    .Z(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5531_ (.A1(\mod.registers.r5[6] ),
    .A2(_2405_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5532_ (.A1(_2411_),
    .A2(_2404_),
    .B(_2412_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5533_ (.I(_2235_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5534_ (.I(_2413_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5535_ (.A1(\mod.registers.r5[7] ),
    .A2(_2405_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5536_ (.A1(_2414_),
    .A2(_2404_),
    .B(_2415_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5537_ (.I(_2244_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5538_ (.I(_2416_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5539_ (.I(_2388_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5540_ (.I(_2390_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5541_ (.A1(\mod.registers.r5[8] ),
    .A2(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5542_ (.A1(_2417_),
    .A2(_2418_),
    .B(_2420_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5543_ (.I(_2253_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5544_ (.I(_2421_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5545_ (.A1(\mod.registers.r5[9] ),
    .A2(_2419_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5546_ (.A1(_2422_),
    .A2(_2418_),
    .B(_2423_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5547_ (.I(_2260_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5548_ (.I(_2424_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5549_ (.A1(\mod.registers.r5[10] ),
    .A2(_2419_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5550_ (.A1(_2425_),
    .A2(_2418_),
    .B(_2426_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5551_ (.I(_2267_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5552_ (.I(_2427_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5553_ (.A1(\mod.registers.r5[11] ),
    .A2(_2419_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5554_ (.A1(_2428_),
    .A2(_2418_),
    .B(_2429_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5555_ (.I(_2275_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5556_ (.I(_2430_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5557_ (.I(_2388_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5558_ (.I(_2390_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5559_ (.A1(\mod.registers.r5[12] ),
    .A2(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5560_ (.A1(_2431_),
    .A2(_2432_),
    .B(_2434_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5561_ (.I(_2283_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5562_ (.I(_2435_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5563_ (.A1(\mod.registers.r5[13] ),
    .A2(_2433_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5564_ (.A1(_2436_),
    .A2(_2432_),
    .B(_2437_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5565_ (.I(_2289_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5566_ (.I(_2438_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5567_ (.A1(\mod.registers.r5[14] ),
    .A2(_2433_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5568_ (.A1(_2439_),
    .A2(_2432_),
    .B(_2440_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5569_ (.I(_2295_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5570_ (.I(_2441_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5571_ (.A1(\mod.registers.r5[15] ),
    .A2(_2433_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5572_ (.A1(_2442_),
    .A2(_2432_),
    .B(_2443_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5573_ (.A1(_2299_),
    .A2(_2356_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5574_ (.I(_2444_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5575_ (.I(_2445_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5576_ (.I(_2444_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5577_ (.I(_2447_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5578_ (.A1(\mod.registers.r6[0] ),
    .A2(_2448_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5579_ (.A1(_2386_),
    .A2(_2446_),
    .B(_2449_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5580_ (.A1(\mod.registers.r6[1] ),
    .A2(_2448_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5581_ (.A1(_2394_),
    .A2(_2446_),
    .B(_2450_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5582_ (.A1(\mod.registers.r6[2] ),
    .A2(_2448_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5583_ (.A1(_2397_),
    .A2(_2446_),
    .B(_2451_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5584_ (.A1(\mod.registers.r6[3] ),
    .A2(_2448_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5585_ (.A1(_2400_),
    .A2(_2446_),
    .B(_2452_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5586_ (.I(_2445_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5587_ (.I(_2447_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5588_ (.A1(\mod.registers.r6[4] ),
    .A2(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5589_ (.A1(_2403_),
    .A2(_2453_),
    .B(_2455_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5590_ (.A1(\mod.registers.r6[5] ),
    .A2(_2454_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5591_ (.A1(_2408_),
    .A2(_2453_),
    .B(_2456_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5592_ (.A1(\mod.registers.r6[6] ),
    .A2(_2454_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5593_ (.A1(_2411_),
    .A2(_2453_),
    .B(_2457_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5594_ (.A1(\mod.registers.r6[7] ),
    .A2(_2454_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5595_ (.A1(_2414_),
    .A2(_2453_),
    .B(_2458_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5596_ (.I(_2445_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5597_ (.I(_2447_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5598_ (.A1(\mod.registers.r6[8] ),
    .A2(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5599_ (.A1(_2417_),
    .A2(_2459_),
    .B(_2461_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5600_ (.A1(\mod.registers.r6[9] ),
    .A2(_2460_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5601_ (.A1(_2422_),
    .A2(_2459_),
    .B(_2462_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5602_ (.A1(\mod.registers.r6[10] ),
    .A2(_2460_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5603_ (.A1(_2425_),
    .A2(_2459_),
    .B(_2463_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5604_ (.A1(\mod.registers.r6[11] ),
    .A2(_2460_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5605_ (.A1(_2428_),
    .A2(_2459_),
    .B(_2464_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5606_ (.I(_2445_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5607_ (.I(_2447_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5608_ (.A1(\mod.registers.r6[12] ),
    .A2(_2466_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5609_ (.A1(_2431_),
    .A2(_2465_),
    .B(_2467_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5610_ (.A1(\mod.registers.r6[13] ),
    .A2(_2466_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5611_ (.A1(_2436_),
    .A2(_2465_),
    .B(_2468_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5612_ (.A1(\mod.registers.r6[14] ),
    .A2(_2466_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5613_ (.A1(_2439_),
    .A2(_2465_),
    .B(_2469_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5614_ (.A1(\mod.registers.r6[15] ),
    .A2(_2466_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5615_ (.A1(_2442_),
    .A2(_2465_),
    .B(_2470_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5616_ (.A1(_2327_),
    .A2(_2356_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5617_ (.I(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5618_ (.I(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5619_ (.I(_2471_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5620_ (.I(_2474_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5621_ (.A1(\mod.registers.r7[0] ),
    .A2(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5622_ (.A1(_2386_),
    .A2(_2473_),
    .B(_2476_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5623_ (.A1(\mod.registers.r7[1] ),
    .A2(_2475_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5624_ (.A1(_2394_),
    .A2(_2473_),
    .B(_2477_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5625_ (.A1(\mod.registers.r7[2] ),
    .A2(_2475_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5626_ (.A1(_2397_),
    .A2(_2473_),
    .B(_2478_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5627_ (.A1(\mod.registers.r7[3] ),
    .A2(_2475_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5628_ (.A1(_2400_),
    .A2(_2473_),
    .B(_2479_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5629_ (.I(_2472_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5630_ (.I(_2474_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5631_ (.A1(\mod.registers.r7[4] ),
    .A2(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5632_ (.A1(_2403_),
    .A2(_2480_),
    .B(_2482_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5633_ (.A1(\mod.registers.r7[5] ),
    .A2(_2481_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5634_ (.A1(_2408_),
    .A2(_2480_),
    .B(_2483_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5635_ (.A1(\mod.registers.r7[6] ),
    .A2(_2481_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5636_ (.A1(_2411_),
    .A2(_2480_),
    .B(_2484_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5637_ (.A1(\mod.registers.r7[7] ),
    .A2(_2481_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5638_ (.A1(_2414_),
    .A2(_2480_),
    .B(_2485_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5639_ (.I(_2472_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5640_ (.I(_2474_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5641_ (.A1(\mod.registers.r7[8] ),
    .A2(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5642_ (.A1(_2417_),
    .A2(_2486_),
    .B(_2488_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5643_ (.A1(\mod.registers.r7[9] ),
    .A2(_2487_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5644_ (.A1(_2422_),
    .A2(_2486_),
    .B(_2489_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5645_ (.A1(\mod.registers.r7[10] ),
    .A2(_2487_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5646_ (.A1(_2425_),
    .A2(_2486_),
    .B(_2490_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5647_ (.A1(\mod.registers.r7[11] ),
    .A2(_2487_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5648_ (.A1(_2428_),
    .A2(_2486_),
    .B(_2491_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5649_ (.I(_2472_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5650_ (.I(_2474_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5651_ (.A1(\mod.registers.r7[12] ),
    .A2(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5652_ (.A1(_2431_),
    .A2(_2492_),
    .B(_2494_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5653_ (.A1(\mod.registers.r7[13] ),
    .A2(_2493_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5654_ (.A1(_2436_),
    .A2(_2492_),
    .B(_2495_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5655_ (.A1(\mod.registers.r7[14] ),
    .A2(_2493_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5656_ (.A1(_2439_),
    .A2(_2492_),
    .B(_2496_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(\mod.registers.r7[15] ),
    .A2(_2493_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_2442_),
    .A2(_2492_),
    .B(_2497_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5659_ (.I(_2149_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5660_ (.A1(_2146_),
    .A2(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(_2357_),
    .A2(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5662_ (.I(_2500_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5663_ (.I(_2501_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5664_ (.I(_2500_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5665_ (.I(_2503_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5666_ (.A1(\mod.registers.r8[0] ),
    .A2(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5667_ (.A1(_2386_),
    .A2(_2502_),
    .B(_2505_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(\mod.registers.r8[1] ),
    .A2(_2504_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5669_ (.A1(_2394_),
    .A2(_2502_),
    .B(_2506_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5670_ (.A1(\mod.registers.r8[2] ),
    .A2(_2504_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5671_ (.A1(_2397_),
    .A2(_2502_),
    .B(_2507_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5672_ (.A1(\mod.registers.r8[3] ),
    .A2(_2504_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5673_ (.A1(_2400_),
    .A2(_2502_),
    .B(_2508_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5674_ (.I(_2501_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5675_ (.I(_2503_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5676_ (.A1(\mod.registers.r8[4] ),
    .A2(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5677_ (.A1(_2403_),
    .A2(_2509_),
    .B(_2511_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5678_ (.A1(\mod.registers.r8[5] ),
    .A2(_2510_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5679_ (.A1(_2408_),
    .A2(_2509_),
    .B(_2512_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(\mod.registers.r8[6] ),
    .A2(_2510_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5681_ (.A1(_2411_),
    .A2(_2509_),
    .B(_2513_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5682_ (.A1(\mod.registers.r8[7] ),
    .A2(_2510_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5683_ (.A1(_2414_),
    .A2(_2509_),
    .B(_2514_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5684_ (.I(_2501_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5685_ (.I(_2503_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5686_ (.A1(\mod.registers.r8[8] ),
    .A2(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5687_ (.A1(_2417_),
    .A2(_2515_),
    .B(_2517_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(\mod.registers.r8[9] ),
    .A2(_2516_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5689_ (.A1(_2422_),
    .A2(_2515_),
    .B(_2518_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5690_ (.A1(\mod.registers.r8[10] ),
    .A2(_2516_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5691_ (.A1(_2425_),
    .A2(_2515_),
    .B(_2519_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5692_ (.A1(\mod.registers.r8[11] ),
    .A2(_2516_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5693_ (.A1(_2428_),
    .A2(_2515_),
    .B(_2520_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_2501_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5695_ (.I(_2503_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5696_ (.A1(\mod.registers.r8[12] ),
    .A2(_2522_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5697_ (.A1(_2431_),
    .A2(_2521_),
    .B(_2523_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5698_ (.A1(\mod.registers.r8[13] ),
    .A2(_2522_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5699_ (.A1(_2436_),
    .A2(_2521_),
    .B(_2524_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5700_ (.A1(\mod.registers.r8[14] ),
    .A2(_2522_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5701_ (.A1(_2439_),
    .A2(_2521_),
    .B(_2525_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5702_ (.A1(\mod.registers.r8[15] ),
    .A2(_2522_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5703_ (.A1(_2442_),
    .A2(_2521_),
    .B(_2526_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5704_ (.I(_2176_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5705_ (.A1(_2161_),
    .A2(_2499_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5706_ (.I(_2528_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_2529_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5708_ (.I(_2528_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5709_ (.I(_2531_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5710_ (.A1(\mod.registers.r9[0] ),
    .A2(_2532_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5711_ (.A1(_2527_),
    .A2(_2530_),
    .B(_2533_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5712_ (.I(_2185_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5713_ (.A1(\mod.registers.r9[1] ),
    .A2(_2532_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5714_ (.A1(_2534_),
    .A2(_2530_),
    .B(_2535_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_2193_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5716_ (.A1(\mod.registers.r9[2] ),
    .A2(_2532_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5717_ (.A1(_2536_),
    .A2(_2530_),
    .B(_2537_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5718_ (.I(_2198_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5719_ (.A1(\mod.registers.r9[3] ),
    .A2(_2532_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5720_ (.A1(_2538_),
    .A2(_2530_),
    .B(_2539_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5721_ (.I(_2204_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5722_ (.I(_2529_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_2531_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5724_ (.A1(\mod.registers.r9[4] ),
    .A2(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5725_ (.A1(_2540_),
    .A2(_2541_),
    .B(_2543_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5726_ (.I(_2217_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5727_ (.A1(\mod.registers.r9[5] ),
    .A2(_2542_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5728_ (.A1(_2544_),
    .A2(_2541_),
    .B(_2545_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5729_ (.I(_2228_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5730_ (.A1(\mod.registers.r9[6] ),
    .A2(_2542_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5731_ (.A1(_2546_),
    .A2(_2541_),
    .B(_2547_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5732_ (.I(_2235_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5733_ (.A1(\mod.registers.r9[7] ),
    .A2(_2542_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5734_ (.A1(_2548_),
    .A2(_2541_),
    .B(_2549_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5735_ (.I(_2244_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5736_ (.I(_2529_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_2531_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5738_ (.A1(\mod.registers.r9[8] ),
    .A2(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5739_ (.A1(_2550_),
    .A2(_2551_),
    .B(_2553_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5740_ (.I(_2253_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5741_ (.A1(\mod.registers.r9[9] ),
    .A2(_2552_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5742_ (.A1(_2554_),
    .A2(_2551_),
    .B(_2555_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5743_ (.I(_2260_),
    .Z(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(\mod.registers.r9[10] ),
    .A2(_2552_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5745_ (.A1(_2556_),
    .A2(_2551_),
    .B(_2557_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_2267_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5747_ (.A1(\mod.registers.r9[11] ),
    .A2(_2552_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5748_ (.A1(_2558_),
    .A2(_2551_),
    .B(_2559_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5749_ (.I(_2275_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5750_ (.I(_2529_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5751_ (.I(_2531_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5752_ (.A1(\mod.registers.r9[12] ),
    .A2(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5753_ (.A1(_2560_),
    .A2(_2561_),
    .B(_2563_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5754_ (.I(_2283_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5755_ (.A1(\mod.registers.r9[13] ),
    .A2(_2562_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5756_ (.A1(_2564_),
    .A2(_2561_),
    .B(_2565_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5757_ (.I(_2289_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5758_ (.A1(\mod.registers.r9[14] ),
    .A2(_2562_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5759_ (.A1(_2566_),
    .A2(_2561_),
    .B(_2567_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5760_ (.I(_2295_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5761_ (.A1(\mod.registers.r9[15] ),
    .A2(_2562_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5762_ (.A1(_2568_),
    .A2(_2561_),
    .B(_2569_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5763_ (.A1(_2299_),
    .A2(_2499_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5764_ (.I(_2570_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5765_ (.I(_2571_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5766_ (.I(_2570_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5767_ (.I(_2573_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5768_ (.A1(\mod.registers.r10[0] ),
    .A2(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5769_ (.A1(_2527_),
    .A2(_2572_),
    .B(_2575_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5770_ (.A1(\mod.registers.r10[1] ),
    .A2(_2574_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5771_ (.A1(_2534_),
    .A2(_2572_),
    .B(_2576_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5772_ (.A1(\mod.registers.r10[2] ),
    .A2(_2574_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5773_ (.A1(_2536_),
    .A2(_2572_),
    .B(_2577_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5774_ (.A1(\mod.registers.r10[3] ),
    .A2(_2574_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5775_ (.A1(_2538_),
    .A2(_2572_),
    .B(_2578_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5776_ (.I(_2571_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5777_ (.I(_2573_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5778_ (.A1(\mod.registers.r10[4] ),
    .A2(_2580_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5779_ (.A1(_2540_),
    .A2(_2579_),
    .B(_2581_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5780_ (.A1(\mod.registers.r10[5] ),
    .A2(_2580_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5781_ (.A1(_2544_),
    .A2(_2579_),
    .B(_2582_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5782_ (.A1(\mod.registers.r10[6] ),
    .A2(_2580_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5783_ (.A1(_2546_),
    .A2(_2579_),
    .B(_2583_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5784_ (.A1(\mod.registers.r10[7] ),
    .A2(_2580_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5785_ (.A1(_2548_),
    .A2(_2579_),
    .B(_2584_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5786_ (.I(_2571_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5787_ (.I(_2573_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5788_ (.A1(\mod.registers.r10[8] ),
    .A2(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5789_ (.A1(_2550_),
    .A2(_2585_),
    .B(_2587_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5790_ (.A1(\mod.registers.r10[9] ),
    .A2(_2586_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5791_ (.A1(_2554_),
    .A2(_2585_),
    .B(_2588_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5792_ (.A1(\mod.registers.r10[10] ),
    .A2(_2586_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5793_ (.A1(_2556_),
    .A2(_2585_),
    .B(_2589_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5794_ (.A1(\mod.registers.r10[11] ),
    .A2(_2586_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5795_ (.A1(_2558_),
    .A2(_2585_),
    .B(_2590_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5796_ (.I(_2571_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5797_ (.I(_2573_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5798_ (.A1(\mod.registers.r10[12] ),
    .A2(_2592_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5799_ (.A1(_2560_),
    .A2(_2591_),
    .B(_2593_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5800_ (.A1(\mod.registers.r10[13] ),
    .A2(_2592_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5801_ (.A1(_2564_),
    .A2(_2591_),
    .B(_2594_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5802_ (.A1(\mod.registers.r10[14] ),
    .A2(_2592_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5803_ (.A1(_2566_),
    .A2(_2591_),
    .B(_2595_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5804_ (.A1(\mod.registers.r10[15] ),
    .A2(_2592_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5805_ (.A1(_2568_),
    .A2(_2591_),
    .B(_2596_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5806_ (.A1(_2327_),
    .A2(_2499_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5807_ (.I(_2597_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5808_ (.I(_2598_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5809_ (.I(_2597_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5810_ (.I(_2600_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(\mod.registers.r11[0] ),
    .A2(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5812_ (.A1(_2527_),
    .A2(_2599_),
    .B(_2602_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5813_ (.A1(\mod.registers.r11[1] ),
    .A2(_2601_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5814_ (.A1(_2534_),
    .A2(_2599_),
    .B(_2603_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(\mod.registers.r11[2] ),
    .A2(_2601_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5816_ (.A1(_2536_),
    .A2(_2599_),
    .B(_2604_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(\mod.registers.r11[3] ),
    .A2(_2601_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5818_ (.A1(_2538_),
    .A2(_2599_),
    .B(_2605_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5819_ (.I(_2598_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5820_ (.I(_2600_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5821_ (.A1(\mod.registers.r11[4] ),
    .A2(_2607_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5822_ (.A1(_2540_),
    .A2(_2606_),
    .B(_2608_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5823_ (.A1(\mod.registers.r11[5] ),
    .A2(_2607_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5824_ (.A1(_2544_),
    .A2(_2606_),
    .B(_2609_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5825_ (.A1(\mod.registers.r11[6] ),
    .A2(_2607_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5826_ (.A1(_2546_),
    .A2(_2606_),
    .B(_2610_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5827_ (.A1(\mod.registers.r11[7] ),
    .A2(_2607_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5828_ (.A1(_2548_),
    .A2(_2606_),
    .B(_2611_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5829_ (.I(_2598_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5830_ (.I(_2600_),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5831_ (.A1(\mod.registers.r11[8] ),
    .A2(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5832_ (.A1(_2550_),
    .A2(_2612_),
    .B(_2614_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5833_ (.A1(\mod.registers.r11[9] ),
    .A2(_2613_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5834_ (.A1(_2554_),
    .A2(_2612_),
    .B(_2615_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5835_ (.A1(\mod.registers.r11[10] ),
    .A2(_2613_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5836_ (.A1(_2556_),
    .A2(_2612_),
    .B(_2616_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5837_ (.A1(\mod.registers.r11[11] ),
    .A2(_2613_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5838_ (.A1(_2558_),
    .A2(_2612_),
    .B(_2617_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5839_ (.I(_2598_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5840_ (.I(_2600_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5841_ (.A1(\mod.registers.r11[12] ),
    .A2(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5842_ (.A1(_2560_),
    .A2(_2618_),
    .B(_2620_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5843_ (.A1(\mod.registers.r11[13] ),
    .A2(_2619_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5844_ (.A1(_2564_),
    .A2(_2618_),
    .B(_2621_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5845_ (.A1(\mod.registers.r11[14] ),
    .A2(_2619_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5846_ (.A1(_2566_),
    .A2(_2618_),
    .B(_2622_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5847_ (.A1(\mod.registers.r11[15] ),
    .A2(_2619_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5848_ (.A1(_2568_),
    .A2(_2618_),
    .B(_2623_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5849_ (.A1(_2355_),
    .A2(_2498_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5850_ (.A1(_2357_),
    .A2(_2624_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5851_ (.I(_2625_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5852_ (.I(_2626_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5853_ (.I(_2625_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5854_ (.I(_2628_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5855_ (.A1(\mod.registers.r12[0] ),
    .A2(_2629_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5856_ (.A1(_2527_),
    .A2(_2627_),
    .B(_2630_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5857_ (.A1(\mod.registers.r12[1] ),
    .A2(_2629_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5858_ (.A1(_2534_),
    .A2(_2627_),
    .B(_2631_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5859_ (.A1(\mod.registers.r12[2] ),
    .A2(_2629_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5860_ (.A1(_2536_),
    .A2(_2627_),
    .B(_2632_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5861_ (.A1(\mod.registers.r12[3] ),
    .A2(_2629_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5862_ (.A1(_2538_),
    .A2(_2627_),
    .B(_2633_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5863_ (.I(_2626_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5864_ (.I(_2628_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5865_ (.A1(\mod.registers.r12[4] ),
    .A2(_2635_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5866_ (.A1(_2540_),
    .A2(_2634_),
    .B(_2636_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5867_ (.A1(\mod.registers.r12[5] ),
    .A2(_2635_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5868_ (.A1(_2544_),
    .A2(_2634_),
    .B(_2637_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5869_ (.A1(\mod.registers.r12[6] ),
    .A2(_2635_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5870_ (.A1(_2546_),
    .A2(_2634_),
    .B(_2638_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5871_ (.A1(\mod.registers.r12[7] ),
    .A2(_2635_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5872_ (.A1(_2548_),
    .A2(_2634_),
    .B(_2639_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5873_ (.I(_2626_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5874_ (.I(_2628_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5875_ (.A1(\mod.registers.r12[8] ),
    .A2(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5876_ (.A1(_2550_),
    .A2(_2640_),
    .B(_2642_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5877_ (.A1(\mod.registers.r12[9] ),
    .A2(_2641_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5878_ (.A1(_2554_),
    .A2(_2640_),
    .B(_2643_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5879_ (.A1(\mod.registers.r12[10] ),
    .A2(_2641_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5880_ (.A1(_2556_),
    .A2(_2640_),
    .B(_2644_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5881_ (.A1(\mod.registers.r12[11] ),
    .A2(_2641_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5882_ (.A1(_2558_),
    .A2(_2640_),
    .B(_2645_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5883_ (.I(_2626_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5884_ (.I(_2628_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5885_ (.A1(\mod.registers.r12[12] ),
    .A2(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5886_ (.A1(_2560_),
    .A2(_2646_),
    .B(_2648_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5887_ (.A1(\mod.registers.r12[13] ),
    .A2(_2647_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5888_ (.A1(_2564_),
    .A2(_2646_),
    .B(_2649_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5889_ (.A1(\mod.registers.r12[14] ),
    .A2(_2647_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5890_ (.A1(_2566_),
    .A2(_2646_),
    .B(_2650_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(\mod.registers.r12[15] ),
    .A2(_2647_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5892_ (.A1(_2568_),
    .A2(_2646_),
    .B(_2651_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(_2161_),
    .A2(_2624_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5894_ (.I(_2652_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5895_ (.I(_2653_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5896_ (.I(_2652_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5897_ (.I(_2655_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5898_ (.A1(\mod.registers.r13[0] ),
    .A2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5899_ (.A1(_2385_),
    .A2(_2654_),
    .B(_2657_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5900_ (.A1(\mod.registers.r13[1] ),
    .A2(_2656_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5901_ (.A1(_2393_),
    .A2(_2654_),
    .B(_2658_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5902_ (.A1(\mod.registers.r13[2] ),
    .A2(_2656_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5903_ (.A1(_2396_),
    .A2(_2654_),
    .B(_2659_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5904_ (.A1(\mod.registers.r13[3] ),
    .A2(_2656_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5905_ (.A1(_2399_),
    .A2(_2654_),
    .B(_2660_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5906_ (.I(_2653_),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5907_ (.I(_2655_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5908_ (.A1(\mod.registers.r13[4] ),
    .A2(_2662_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5909_ (.A1(_2402_),
    .A2(_2661_),
    .B(_2663_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5910_ (.A1(\mod.registers.r13[5] ),
    .A2(_2662_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5911_ (.A1(_2407_),
    .A2(_2661_),
    .B(_2664_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5912_ (.A1(\mod.registers.r13[6] ),
    .A2(_2662_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5913_ (.A1(_2410_),
    .A2(_2661_),
    .B(_2665_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5914_ (.A1(\mod.registers.r13[7] ),
    .A2(_2662_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5915_ (.A1(_2413_),
    .A2(_2661_),
    .B(_2666_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5916_ (.I(_2653_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5917_ (.I(_2655_),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5918_ (.A1(\mod.registers.r13[8] ),
    .A2(_2668_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5919_ (.A1(_2416_),
    .A2(_2667_),
    .B(_2669_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5920_ (.A1(\mod.registers.r13[9] ),
    .A2(_2668_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5921_ (.A1(_2421_),
    .A2(_2667_),
    .B(_2670_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5922_ (.A1(\mod.registers.r13[10] ),
    .A2(_2668_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5923_ (.A1(_2424_),
    .A2(_2667_),
    .B(_2671_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5924_ (.A1(\mod.registers.r13[11] ),
    .A2(_2668_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5925_ (.A1(_2427_),
    .A2(_2667_),
    .B(_2672_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5926_ (.I(_2653_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5927_ (.I(_2655_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5928_ (.A1(\mod.registers.r13[12] ),
    .A2(_2674_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5929_ (.A1(_2430_),
    .A2(_2673_),
    .B(_2675_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5930_ (.A1(\mod.registers.r13[13] ),
    .A2(_2674_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5931_ (.A1(_2435_),
    .A2(_2673_),
    .B(_2676_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5932_ (.A1(\mod.registers.r13[14] ),
    .A2(_2674_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5933_ (.A1(_2438_),
    .A2(_2673_),
    .B(_2677_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5934_ (.A1(\mod.registers.r13[15] ),
    .A2(_2674_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5935_ (.A1(_2441_),
    .A2(_2673_),
    .B(_2678_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5936_ (.A1(_2299_),
    .A2(_2624_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5937_ (.I(_2679_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5938_ (.I(_2680_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5939_ (.I(_2679_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5940_ (.I(_2682_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5941_ (.A1(\mod.registers.r14[0] ),
    .A2(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5942_ (.A1(_2385_),
    .A2(_2681_),
    .B(_2684_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5943_ (.A1(\mod.registers.r14[1] ),
    .A2(_2683_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5944_ (.A1(_2393_),
    .A2(_2681_),
    .B(_2685_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5945_ (.A1(\mod.registers.r14[2] ),
    .A2(_2683_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5946_ (.A1(_2396_),
    .A2(_2681_),
    .B(_2686_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5947_ (.A1(\mod.registers.r14[3] ),
    .A2(_2683_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5948_ (.A1(_2399_),
    .A2(_2681_),
    .B(_2687_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5949_ (.I(_2680_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_2682_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5951_ (.A1(\mod.registers.r14[4] ),
    .A2(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5952_ (.A1(_2402_),
    .A2(_2688_),
    .B(_2690_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5953_ (.A1(\mod.registers.r14[5] ),
    .A2(_2689_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5954_ (.A1(_2407_),
    .A2(_2688_),
    .B(_2691_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5955_ (.A1(\mod.registers.r14[6] ),
    .A2(_2689_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5956_ (.A1(_2410_),
    .A2(_2688_),
    .B(_2692_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5957_ (.A1(\mod.registers.r14[7] ),
    .A2(_2689_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5958_ (.A1(_2413_),
    .A2(_2688_),
    .B(_2693_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5959_ (.I(_2680_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_2682_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5961_ (.A1(\mod.registers.r14[8] ),
    .A2(_2695_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5962_ (.A1(_2416_),
    .A2(_2694_),
    .B(_2696_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5963_ (.A1(\mod.registers.r14[9] ),
    .A2(_2695_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5964_ (.A1(_2421_),
    .A2(_2694_),
    .B(_2697_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5965_ (.A1(\mod.registers.r14[10] ),
    .A2(_2695_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5966_ (.A1(_2424_),
    .A2(_2694_),
    .B(_2698_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5967_ (.A1(\mod.registers.r14[11] ),
    .A2(_2695_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5968_ (.A1(_2427_),
    .A2(_2694_),
    .B(_2699_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5969_ (.I(_2680_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5970_ (.I(_2682_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5971_ (.A1(\mod.registers.r14[12] ),
    .A2(_2701_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5972_ (.A1(_2430_),
    .A2(_2700_),
    .B(_2702_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5973_ (.A1(\mod.registers.r14[13] ),
    .A2(_2701_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5974_ (.A1(_2435_),
    .A2(_2700_),
    .B(_2703_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5975_ (.A1(\mod.registers.r14[14] ),
    .A2(_2701_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5976_ (.A1(_2438_),
    .A2(_2700_),
    .B(_2704_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5977_ (.A1(\mod.registers.r14[15] ),
    .A2(_2701_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5978_ (.A1(_2441_),
    .A2(_2700_),
    .B(_2705_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5979_ (.I(net11),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5980_ (.I(_2706_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5981_ (.I(_2707_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5982_ (.I(_2708_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5983_ (.I(_2708_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5984_ (.I(_2708_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5985_ (.A1(_1895_),
    .A2(_1884_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5986_ (.A1(\mod.valid0 ),
    .A2(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5987_ (.I(net12),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5988_ (.A1(_2711_),
    .A2(_1884_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5989_ (.I(_2712_),
    .Z(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5990_ (.I(_2713_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5991_ (.I(_2706_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_2715_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5993_ (.A1(_2710_),
    .A2(_2714_),
    .B(_2716_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5994_ (.A1(\mod.valid0 ),
    .A2(_2709_),
    .A3(_2151_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5995_ (.I(_2717_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_2718_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5997_ (.I(_2712_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5998_ (.A1(\mod.valid1 ),
    .A2(_2709_),
    .A3(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5999_ (.A1(_2719_),
    .A2(_2721_),
    .B(_2716_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_2711_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_2722_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6002_ (.A1(_2723_),
    .A2(\mod.pc0[0] ),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6003_ (.I(_2711_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6004_ (.I(_2725_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6005_ (.A1(_2726_),
    .A2(_1903_),
    .B(_0003_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6006_ (.A1(_2724_),
    .A2(_2727_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6007_ (.I(_2711_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6008_ (.I(_2728_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6009_ (.I(_2729_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6010_ (.I(_2140_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6011_ (.A1(_2723_),
    .A2(\mod.pc0[1] ),
    .B(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6012_ (.A1(_2730_),
    .A2(_1928_),
    .B(_2732_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6013_ (.A1(_2726_),
    .A2(_1947_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_2728_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6015_ (.A1(_2734_),
    .A2(\mod.pc0[2] ),
    .B(_2731_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6016_ (.A1(_2733_),
    .A2(_2735_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6017_ (.I(_2728_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6018_ (.A1(_2736_),
    .A2(_1959_),
    .A3(_1965_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6019_ (.A1(_2734_),
    .A2(\mod.pc0[3] ),
    .B(_2737_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6020_ (.A1(_2708_),
    .A2(_2738_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6021_ (.A1(_2723_),
    .A2(\mod.pc0[4] ),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6022_ (.A1(_2726_),
    .A2(_1983_),
    .B(_2731_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6023_ (.A1(_2739_),
    .A2(_2740_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6024_ (.I(_2706_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6025_ (.I(_2741_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6026_ (.I(_2742_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6027_ (.A1(_2736_),
    .A2(_1998_),
    .A3(_2001_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6028_ (.A1(_2734_),
    .A2(\mod.pc0[5] ),
    .B(_2744_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6029_ (.A1(_2743_),
    .A2(_2745_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6030_ (.I(_2722_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6031_ (.A1(_2736_),
    .A2(_2016_),
    .A3(_2019_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6032_ (.A1(_2746_),
    .A2(\mod.pc0[6] ),
    .B(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6033_ (.A1(_2743_),
    .A2(_2748_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6034_ (.A1(_2736_),
    .A2(_2032_),
    .A3(_2035_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6035_ (.A1(_2746_),
    .A2(\mod.pc0[7] ),
    .B(_2749_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6036_ (.A1(_2743_),
    .A2(_2750_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6037_ (.A1(_2729_),
    .A2(\mod.pc0[8] ),
    .B(_2731_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6038_ (.A1(_2730_),
    .A2(_2053_),
    .B(_2751_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6039_ (.I(_2139_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6040_ (.I(_2752_),
    .Z(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6041_ (.I(_2753_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6042_ (.A1(_2729_),
    .A2(\mod.pc0[9] ),
    .B(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6043_ (.A1(_2730_),
    .A2(_2069_),
    .B(_2755_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6044_ (.A1(_2722_),
    .A2(_2084_),
    .A3(_2087_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6045_ (.A1(_2746_),
    .A2(\mod.pc0[10] ),
    .B(_2756_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6046_ (.A1(_2743_),
    .A2(_2757_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6047_ (.A1(_2729_),
    .A2(\mod.pc0[11] ),
    .B(_2754_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6048_ (.A1(_2730_),
    .A2(_2105_),
    .B(_2758_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6049_ (.I(_2741_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6050_ (.I(_2759_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6051_ (.A1(_2722_),
    .A2(_2114_),
    .A3(_2117_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6052_ (.A1(_2746_),
    .A2(\mod.pc0[12] ),
    .B(_2761_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6053_ (.A1(_2760_),
    .A2(_2762_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6054_ (.A1(\mod.pc0[13] ),
    .A2(_2723_),
    .B(_2754_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6055_ (.A1(_2734_),
    .A2(_2134_),
    .B(_2763_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6056_ (.A1(_2725_),
    .A2(_1899_),
    .Z(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6057_ (.I(_2764_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6058_ (.I(_2765_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6059_ (.I(_2764_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6060_ (.I(_1389_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6061_ (.I(_1788_),
    .Z(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6062_ (.A1(_2768_),
    .A2(_2769_),
    .B(\mod.pc[0] ),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6063_ (.A1(_1797_),
    .A2(_2770_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6064_ (.A1(_2767_),
    .A2(_2771_),
    .B(_2754_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6065_ (.A1(_1893_),
    .A2(_2766_),
    .B(_2772_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6066_ (.A1(_2726_),
    .A2(_1900_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6067_ (.I(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6068_ (.A1(_1911_),
    .A2(_2004_),
    .A3(_1920_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6069_ (.A1(_1926_),
    .A2(_2775_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6070_ (.A1(_2771_),
    .A2(_2776_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6071_ (.I(_2753_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6072_ (.A1(\mod.pc[1] ),
    .A2(_2774_),
    .B(_2778_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6073_ (.A1(_2774_),
    .A2(_2777_),
    .B(_2779_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6074_ (.I(_2765_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6075_ (.I(\mod.pc[1] ),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6076_ (.A1(_2781_),
    .A2(_1913_),
    .B1(_1797_),
    .B2(_2770_),
    .C(_2775_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6077_ (.I(_2782_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6078_ (.A1(_2768_),
    .A2(_2004_),
    .B(\mod.pc[2] ),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6079_ (.A1(_1943_),
    .A2(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6080_ (.A1(_2783_),
    .A2(_2785_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6081_ (.A1(_2765_),
    .A2(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6082_ (.I(_2706_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6083_ (.I(_2788_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6084_ (.A1(_1944_),
    .A2(_2780_),
    .B(_2787_),
    .C(_2789_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6085_ (.A1(_2768_),
    .A2(_2769_),
    .B(\mod.pc[3] ),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6086_ (.A1(_1943_),
    .A2(_2784_),
    .B1(_1959_),
    .B2(_2790_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6087_ (.A1(_2782_),
    .A2(_2791_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6088_ (.A1(_1959_),
    .A2(_2790_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6089_ (.A1(_2783_),
    .A2(_2785_),
    .B(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6090_ (.A1(_2792_),
    .A2(_2794_),
    .B(_2773_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6091_ (.A1(_0003_),
    .A2(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6092_ (.A1(_1962_),
    .A2(_2766_),
    .B(_2796_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6093_ (.A1(_2768_),
    .A2(_2769_),
    .B(\mod.pc[4] ),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6094_ (.A1(_1979_),
    .A2(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6095_ (.A1(_2792_),
    .A2(_2798_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6096_ (.A1(_2767_),
    .A2(_2799_),
    .B(_2778_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6097_ (.A1(_1980_),
    .A2(_2766_),
    .B(_2800_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6098_ (.A1(_2783_),
    .A2(_2791_),
    .A3(_2798_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6099_ (.I(_1389_),
    .Z(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6100_ (.A1(_2802_),
    .A2(_2769_),
    .B(\mod.pc[5] ),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6101_ (.A1(_1998_),
    .A2(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6102_ (.A1(_2801_),
    .A2(_2804_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6103_ (.A1(_2767_),
    .A2(_2805_),
    .B(_2778_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6104_ (.A1(_1999_),
    .A2(_2766_),
    .B(_2806_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6105_ (.A1(_1979_),
    .A2(_2797_),
    .B1(_1998_),
    .B2(_2803_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6106_ (.A1(_2783_),
    .A2(_2791_),
    .A3(_2807_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6107_ (.A1(_2802_),
    .A2(_1885_),
    .B(\mod.pc[6] ),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6108_ (.A1(_2016_),
    .A2(_2809_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6109_ (.A1(_2808_),
    .A2(_2810_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6110_ (.A1(_2767_),
    .A2(_2811_),
    .B(_2778_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6111_ (.A1(_2017_),
    .A2(_2780_),
    .B(_2812_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6112_ (.A1(_2802_),
    .A2(_1885_),
    .B(\mod.pc[7] ),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6113_ (.A1(_2808_),
    .A2(_2810_),
    .B(_2032_),
    .C(_2813_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6114_ (.A1(_2016_),
    .A2(_2809_),
    .B1(_2032_),
    .B2(_2813_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6115_ (.A1(_2782_),
    .A2(_2791_),
    .A3(_2807_),
    .A4(_2815_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6116_ (.I(_2816_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6117_ (.I(_2764_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6118_ (.A1(_2814_),
    .A2(_2817_),
    .B(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6119_ (.A1(_2033_),
    .A2(_2780_),
    .B(_2819_),
    .C(_2789_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6120_ (.A1(_1925_),
    .A2(_2048_),
    .B(_2051_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6121_ (.A1(_2816_),
    .A2(_2820_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6122_ (.I(_2753_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6123_ (.A1(_2765_),
    .A2(_2821_),
    .B(_2822_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6124_ (.A1(_2050_),
    .A2(_2780_),
    .B(_2823_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6125_ (.I(_2818_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6126_ (.A1(\mod.pc[9] ),
    .A2(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6127_ (.A1(_2817_),
    .A2(_2820_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6128_ (.I0(\mod.pc[9] ),
    .I1(_2065_),
    .S(_1894_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6129_ (.I0(\mod.pc[8] ),
    .I1(_2048_),
    .S(_1894_),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6130_ (.A1(_2828_),
    .A2(_2827_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6131_ (.A1(_2826_),
    .A2(_2827_),
    .B1(_2829_),
    .B2(_2817_),
    .C(_2773_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6132_ (.I(_2707_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6133_ (.A1(_2825_),
    .A2(_2830_),
    .B(_2831_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6134_ (.A1(\mod.pc[10] ),
    .A2(_2824_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6135_ (.I(_2816_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6136_ (.A1(_2833_),
    .A2(_2829_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6137_ (.A1(_2802_),
    .A2(_1885_),
    .B(\mod.pc[10] ),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6138_ (.A1(_1913_),
    .A2(_2083_),
    .B(_2835_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6139_ (.A1(_2828_),
    .A2(_2827_),
    .A3(_2836_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6140_ (.I(_2837_),
    .Z(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6141_ (.A1(_2834_),
    .A2(_2836_),
    .B1(_2838_),
    .B2(_2817_),
    .C(_2773_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6142_ (.A1(_2832_),
    .A2(_2839_),
    .B(_2831_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(\mod.pc[11] ),
    .A2(_1914_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6144_ (.A1(_2101_),
    .A2(_2840_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6145_ (.A1(_2833_),
    .A2(_2838_),
    .A3(_2841_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6146_ (.A1(_2833_),
    .A2(_2838_),
    .B(_2841_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6147_ (.A1(_2842_),
    .A2(_2843_),
    .B(_2818_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6148_ (.A1(_2102_),
    .A2(_2824_),
    .B(_2844_),
    .C(_2789_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6149_ (.A1(_2816_),
    .A2(_2837_),
    .A3(_2841_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6150_ (.A1(\mod.pc[12] ),
    .A2(_1914_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6151_ (.A1(_2114_),
    .A2(_2846_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6152_ (.A1(_2845_),
    .A2(_2847_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6153_ (.A1(\mod.pc[12] ),
    .A2(_2774_),
    .B(_2822_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6154_ (.A1(_2774_),
    .A2(_2848_),
    .B(_2849_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6155_ (.A1(_2833_),
    .A2(_2838_),
    .A3(_2841_),
    .A4(_2847_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6156_ (.I(_2130_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6157_ (.A1(_2851_),
    .A2(_2132_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6158_ (.A1(_2850_),
    .A2(_2852_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6159_ (.A1(_2850_),
    .A2(_2852_),
    .B(_2818_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6160_ (.I(_2788_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6161_ (.A1(_2131_),
    .A2(_2824_),
    .B1(_2853_),
    .B2(_2854_),
    .C(_2855_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6162_ (.I(_2151_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(_2856_),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6164_ (.I(_2857_),
    .Z(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6165_ (.I(_2858_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6166_ (.I(_2856_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6167_ (.I(_2860_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6168_ (.A1(\mod.pc_1[0] ),
    .A2(_2861_),
    .B(_2822_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6169_ (.A1(_1893_),
    .A2(_2859_),
    .B(_2862_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6170_ (.A1(\mod.pc_1[1] ),
    .A2(_2861_),
    .B(_2822_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6171_ (.A1(_2781_),
    .A2(_2859_),
    .B(_2863_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6172_ (.I(_2753_),
    .Z(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6173_ (.A1(\mod.pc_1[2] ),
    .A2(_2861_),
    .B(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6174_ (.A1(_1944_),
    .A2(_2859_),
    .B(_2865_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6175_ (.A1(\mod.pc_1[3] ),
    .A2(_2861_),
    .B(_2864_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6176_ (.A1(_1962_),
    .A2(_2859_),
    .B(_2866_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6177_ (.I(_2857_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6178_ (.I(_2867_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6179_ (.I(_2860_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6180_ (.A1(\mod.pc_1[4] ),
    .A2(_2869_),
    .B(_2864_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6181_ (.A1(_1980_),
    .A2(_2868_),
    .B(_2870_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6182_ (.A1(\mod.pc_1[5] ),
    .A2(_2869_),
    .B(_2864_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6183_ (.A1(_1999_),
    .A2(_2868_),
    .B(_2871_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6184_ (.I(_2752_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6185_ (.I(_2872_),
    .Z(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6186_ (.A1(\mod.pc_1[6] ),
    .A2(_2869_),
    .B(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6187_ (.A1(_2017_),
    .A2(_2868_),
    .B(_2874_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6188_ (.A1(\mod.pc_1[7] ),
    .A2(_2869_),
    .B(_2873_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6189_ (.A1(_2033_),
    .A2(_2868_),
    .B(_2875_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6190_ (.I(_2867_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6191_ (.I(_2857_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6192_ (.A1(\mod.pc_1[8] ),
    .A2(_2877_),
    .B(_2873_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6193_ (.A1(_2050_),
    .A2(_2876_),
    .B(_2878_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6194_ (.A1(\mod.pc_1[9] ),
    .A2(_2877_),
    .B(_2873_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6195_ (.A1(_2066_),
    .A2(_2876_),
    .B(_2879_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6196_ (.I(_2872_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6197_ (.A1(\mod.pc_1[10] ),
    .A2(_2877_),
    .B(_2880_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6198_ (.A1(_2085_),
    .A2(_2876_),
    .B(_2881_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6199_ (.A1(\mod.pc_1[11] ),
    .A2(_2877_),
    .B(_2880_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6200_ (.A1(_2102_),
    .A2(_2876_),
    .B(_2882_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6201_ (.I(_2867_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_2857_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6203_ (.A1(\mod.pc_1[12] ),
    .A2(_2884_),
    .B(_2880_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6204_ (.A1(_2115_),
    .A2(_2883_),
    .B(_2885_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6205_ (.A1(\mod.pc_1[13] ),
    .A2(_2884_),
    .B(_2880_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6206_ (.A1(_2131_),
    .A2(_2883_),
    .B(_2886_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6207_ (.I(\mod.instr[0] ),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6208_ (.I(_2717_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6209_ (.I(_2888_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6210_ (.A1(\mod.des.des_dout[0] ),
    .A2(_2889_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6211_ (.I(net13),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6212_ (.I(_2891_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6213_ (.A1(_2887_),
    .A2(_2719_),
    .B1(_2890_),
    .B2(_2892_),
    .C(_2855_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6214_ (.I(\mod.instr[1] ),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6215_ (.A1(\mod.des.des_dout[1] ),
    .A2(_2889_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6216_ (.A1(_2893_),
    .A2(_2719_),
    .B1(_2894_),
    .B2(_2892_),
    .C(_2855_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6217_ (.I(\mod.instr[2] ),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6218_ (.I(_2888_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6219_ (.A1(\mod.des.des_dout[2] ),
    .A2(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6220_ (.I(_2788_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6221_ (.A1(_2895_),
    .A2(_2719_),
    .B1(_2897_),
    .B2(_2892_),
    .C(_2898_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6222_ (.I(\mod.instr[3] ),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6223_ (.I(_2717_),
    .Z(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6224_ (.I(_2900_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6225_ (.A1(\mod.des.des_dout[3] ),
    .A2(_2896_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6226_ (.A1(_2899_),
    .A2(_2901_),
    .B1(_2902_),
    .B2(_2892_),
    .C(_2898_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6227_ (.I(\mod.instr[4] ),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6228_ (.A1(\mod.des.des_dout[4] ),
    .A2(_2896_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6229_ (.I(_2891_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6230_ (.A1(_2903_),
    .A2(_2901_),
    .B1(_2904_),
    .B2(_2905_),
    .C(_2898_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6231_ (.I(\mod.instr[5] ),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6232_ (.A1(\mod.des.des_dout[5] ),
    .A2(_2896_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6233_ (.A1(_2906_),
    .A2(_2901_),
    .B1(_2907_),
    .B2(_2905_),
    .C(_2898_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6234_ (.I(\mod.instr[6] ),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6235_ (.I(_2888_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6236_ (.A1(\mod.des.des_dout[6] ),
    .A2(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6237_ (.I(_2788_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6238_ (.A1(_2908_),
    .A2(_2901_),
    .B1(_2910_),
    .B2(_2905_),
    .C(_2911_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6239_ (.I(\mod.instr[7] ),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6240_ (.I(_2718_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6241_ (.A1(\mod.des.des_dout[7] ),
    .A2(_2909_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6242_ (.A1(_2912_),
    .A2(_2913_),
    .B1(_2914_),
    .B2(_2905_),
    .C(_2911_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6243_ (.I(\mod.instr[8] ),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6244_ (.A1(\mod.des.des_dout[8] ),
    .A2(_2909_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6245_ (.I(_2891_),
    .Z(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6246_ (.A1(_2915_),
    .A2(_2913_),
    .B1(_2916_),
    .B2(_2917_),
    .C(_2911_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6247_ (.I(\mod.instr[9] ),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6248_ (.A1(\mod.des.des_dout[9] ),
    .A2(_2909_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6249_ (.A1(_2918_),
    .A2(_2913_),
    .B1(_2919_),
    .B2(_2917_),
    .C(_2911_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6250_ (.I(\mod.instr[10] ),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6251_ (.I(_2888_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6252_ (.A1(\mod.des.des_dout[10] ),
    .A2(_2921_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6253_ (.I(_2741_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6254_ (.A1(_2920_),
    .A2(_2913_),
    .B1(_2922_),
    .B2(_2917_),
    .C(_2923_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6255_ (.I(\mod.instr[11] ),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6256_ (.I(_2718_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6257_ (.A1(\mod.des.des_dout[11] ),
    .A2(_2921_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6258_ (.A1(_2924_),
    .A2(_2925_),
    .B1(_2926_),
    .B2(_2917_),
    .C(_2923_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6259_ (.I(\mod.instr[12] ),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6260_ (.A1(\mod.des.des_dout[12] ),
    .A2(_2921_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(net13),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6262_ (.A1(_2927_),
    .A2(_2925_),
    .B1(_2928_),
    .B2(_2929_),
    .C(_2923_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6263_ (.I(\mod.instr[13] ),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6264_ (.A1(\mod.des.des_dout[13] ),
    .A2(_2921_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6265_ (.A1(_2930_),
    .A2(_2925_),
    .B1(_2931_),
    .B2(_2929_),
    .C(_2923_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6266_ (.I(\mod.instr[14] ),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6267_ (.I(_2717_),
    .Z(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6268_ (.A1(\mod.des.des_dout[14] ),
    .A2(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6269_ (.I(_2741_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6270_ (.A1(_2932_),
    .A2(_2925_),
    .B1(_2934_),
    .B2(_2929_),
    .C(_2935_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6271_ (.I(\mod.instr[15] ),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6272_ (.I(_2718_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6273_ (.A1(\mod.des.des_dout[15] ),
    .A2(_2933_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6274_ (.A1(_2936_),
    .A2(_2937_),
    .B1(_2938_),
    .B2(_2929_),
    .C(_2935_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6275_ (.I(\mod.instr[16] ),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6276_ (.A1(\mod.des.des_dout[16] ),
    .A2(_2933_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6277_ (.I(net13),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6278_ (.A1(_2939_),
    .A2(_2937_),
    .B1(_2940_),
    .B2(_2941_),
    .C(_2935_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6279_ (.I(\mod.instr[17] ),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6280_ (.A1(\mod.des.des_dout[17] ),
    .A2(_2933_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6281_ (.A1(_2942_),
    .A2(_2937_),
    .B1(_2943_),
    .B2(_2941_),
    .C(_2935_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6282_ (.I(\mod.instr[18] ),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6283_ (.A1(\mod.des.des_dout[18] ),
    .A2(_2900_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6284_ (.A1(_2944_),
    .A2(_2937_),
    .B1(_2945_),
    .B2(_2941_),
    .C(_2742_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6285_ (.I(\mod.instr[19] ),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6286_ (.A1(\mod.des.des_dout[19] ),
    .A2(_2900_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6287_ (.A1(_2946_),
    .A2(_2889_),
    .B1(_2947_),
    .B2(_2941_),
    .C(_2742_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6288_ (.I(\mod.instr[20] ),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6289_ (.A1(\mod.des.des_dout[20] ),
    .A2(_2900_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6290_ (.A1(_2948_),
    .A2(_2889_),
    .B1(_2949_),
    .B2(_2891_),
    .C(_2742_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6291_ (.A1(\mod.valid1 ),
    .A2(_2709_),
    .A3(_2151_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6292_ (.I(_2950_),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6293_ (.I(_2712_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6294_ (.I(_2952_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6295_ (.A1(_1886_),
    .A2(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6296_ (.A1(_2951_),
    .A2(_2954_),
    .B(_2831_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6297_ (.I(_2856_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6298_ (.I(_2955_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6299_ (.A1(_0905_),
    .A2(_2956_),
    .B1(_2951_),
    .B2(\mod.instr[0] ),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6300_ (.A1(_2760_),
    .A2(_2957_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6301_ (.I(_2955_),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6302_ (.A1(_1792_),
    .A2(_2958_),
    .B1(_2951_),
    .B2(\mod.instr[1] ),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6303_ (.A1(_2760_),
    .A2(_2959_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6304_ (.A1(_0903_),
    .A2(_2958_),
    .B1(_2951_),
    .B2(\mod.instr[2] ),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6305_ (.A1(_2760_),
    .A2(_2960_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6306_ (.I(_2759_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6307_ (.I(_2950_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6308_ (.I(_2962_),
    .Z(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6309_ (.A1(\mod.instr_2[3] ),
    .A2(_2958_),
    .B1(_2963_),
    .B2(\mod.instr[3] ),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6310_ (.A1(_2961_),
    .A2(_2964_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6311_ (.A1(\mod.instr_2[4] ),
    .A2(_2958_),
    .B1(_2963_),
    .B2(\mod.instr[4] ),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6312_ (.A1(_2961_),
    .A2(_2965_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6313_ (.I(_1861_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6314_ (.I(_2966_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6315_ (.I(_2955_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6316_ (.A1(_2967_),
    .A2(_2968_),
    .B1(_2963_),
    .B2(\mod.instr[5] ),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6317_ (.A1(_2961_),
    .A2(_2969_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6318_ (.A1(\mod.instr_2[6] ),
    .A2(_2968_),
    .B1(_2963_),
    .B2(\mod.instr[6] ),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6319_ (.A1(_2961_),
    .A2(_2970_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6320_ (.I(_2759_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6321_ (.I(_2962_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6322_ (.A1(_1392_),
    .A2(_2968_),
    .B1(_2972_),
    .B2(\mod.instr[7] ),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6323_ (.A1(_2971_),
    .A2(_2973_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6324_ (.A1(_1391_),
    .A2(_2968_),
    .B1(_2972_),
    .B2(\mod.instr[8] ),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6325_ (.A1(_2971_),
    .A2(_2974_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6326_ (.I(_2955_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6327_ (.A1(_1781_),
    .A2(_2975_),
    .B1(_2972_),
    .B2(\mod.instr[9] ),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6328_ (.A1(_2971_),
    .A2(_2976_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6329_ (.A1(_1805_),
    .A2(_2975_),
    .B1(_2972_),
    .B2(\mod.instr[10] ),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6330_ (.A1(_2971_),
    .A2(_2977_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6331_ (.I(_2759_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6332_ (.I(_2950_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6333_ (.A1(_1808_),
    .A2(_2975_),
    .B1(_2979_),
    .B2(\mod.instr[11] ),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6334_ (.A1(_2978_),
    .A2(_2980_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6335_ (.A1(_0636_),
    .A2(_2975_),
    .B1(_2979_),
    .B2(\mod.instr[12] ),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6336_ (.A1(_2978_),
    .A2(_2981_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6337_ (.I(_2860_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6338_ (.A1(_0846_),
    .A2(_2982_),
    .B1(_2979_),
    .B2(\mod.instr[13] ),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6339_ (.A1(_2978_),
    .A2(_2983_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6340_ (.A1(_1136_),
    .A2(_2982_),
    .B1(_2979_),
    .B2(\mod.instr[14] ),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6341_ (.A1(_2978_),
    .A2(_2984_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6342_ (.I(_2707_),
    .Z(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6343_ (.I(_2950_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6344_ (.A1(_0480_),
    .A2(_2982_),
    .B1(_2986_),
    .B2(\mod.instr[15] ),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6345_ (.A1(_2985_),
    .A2(_2987_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6346_ (.A1(_0616_),
    .A2(_2982_),
    .B1(_2986_),
    .B2(\mod.instr[16] ),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6347_ (.A1(_2985_),
    .A2(_2988_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6348_ (.I(_2860_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6349_ (.A1(_0711_),
    .A2(_2989_),
    .B1(_2986_),
    .B2(\mod.instr[17] ),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6350_ (.A1(_2985_),
    .A2(_2990_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6351_ (.A1(\mod.funct7[0] ),
    .A2(_2989_),
    .B1(_2986_),
    .B2(\mod.instr[18] ),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6352_ (.A1(_2985_),
    .A2(_2991_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6353_ (.I(_2707_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6354_ (.A1(\mod.funct7[1] ),
    .A2(_2989_),
    .B1(_2962_),
    .B2(\mod.instr[19] ),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6355_ (.A1(_2992_),
    .A2(_2993_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6356_ (.A1(_0955_),
    .A2(_2989_),
    .B1(_2962_),
    .B2(\mod.instr[20] ),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6357_ (.A1(_2992_),
    .A2(_2994_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6358_ (.I(_2952_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6359_ (.I(_2872_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6360_ (.A1(\mod.pc_1[0] ),
    .A2(_2995_),
    .B(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6361_ (.A1(_3263_),
    .A2(_2714_),
    .B(_2997_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6362_ (.A1(\mod.pc_1[1] ),
    .A2(_2995_),
    .B(_2996_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6363_ (.A1(_0669_),
    .A2(_2714_),
    .B(_2998_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6364_ (.A1(\mod.pc_1[2] ),
    .A2(_2995_),
    .B(_2996_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6365_ (.A1(_0628_),
    .A2(_2714_),
    .B(_2999_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6366_ (.I(_2713_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6367_ (.I(_2952_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6368_ (.A1(\mod.pc_1[3] ),
    .A2(_3001_),
    .B(_2996_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6369_ (.A1(_0651_),
    .A2(_3000_),
    .B(_3002_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6370_ (.I(_1971_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6371_ (.I(_2872_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6372_ (.A1(\mod.pc_1[4] ),
    .A2(_3001_),
    .B(_3004_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6373_ (.A1(_3003_),
    .A2(_3000_),
    .B(_3005_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6374_ (.A1(\mod.pc_1[5] ),
    .A2(_3001_),
    .B(_3004_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6375_ (.A1(_0580_),
    .A2(_3000_),
    .B(_3006_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6376_ (.I(_2008_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6377_ (.A1(\mod.pc_1[6] ),
    .A2(_3001_),
    .B(_3004_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6378_ (.A1(_3007_),
    .A2(_3000_),
    .B(_3008_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6379_ (.I(_2713_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6380_ (.I(_2952_),
    .Z(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6381_ (.A1(\mod.pc_1[7] ),
    .A2(_3010_),
    .B(_3004_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6382_ (.A1(_0530_),
    .A2(_3009_),
    .B(_3011_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6383_ (.I(_2752_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6384_ (.A1(\mod.pc_1[8] ),
    .A2(_3010_),
    .B(_3012_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6385_ (.A1(_0843_),
    .A2(_3009_),
    .B(_3013_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6386_ (.A1(\mod.pc_1[9] ),
    .A2(_3010_),
    .B(_3012_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6387_ (.A1(_0862_),
    .A2(_3009_),
    .B(_3014_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6388_ (.A1(\mod.pc_1[10] ),
    .A2(_3010_),
    .B(_3012_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6389_ (.A1(_2075_),
    .A2(_3009_),
    .B(_3015_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6390_ (.A1(\mod.pc_1[11] ),
    .A2(_2720_),
    .B(_3012_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6391_ (.A1(_2095_),
    .A2(_2953_),
    .B(_3016_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6392_ (.I(_2752_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6393_ (.A1(\mod.pc_1[12] ),
    .A2(_2720_),
    .B(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6394_ (.A1(_2123_),
    .A2(_2953_),
    .B(_3018_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6395_ (.A1(\mod.pc_1[13] ),
    .A2(_2720_),
    .B(_3017_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6396_ (.A1(_0758_),
    .A2(_2953_),
    .B(_3019_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6397_ (.A1(\mod.valid_out3 ),
    .A2(_2153_),
    .A3(_2713_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6398_ (.A1(_2152_),
    .A2(_3020_),
    .B(_2831_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6399_ (.A1(net20),
    .A2(_2152_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6400_ (.A1(_1886_),
    .A2(_1798_),
    .A3(_3249_),
    .A4(_2858_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6401_ (.I(_2715_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6402_ (.A1(_3021_),
    .A2(_3022_),
    .B(_3023_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6403_ (.A1(\mod.ri_3 ),
    .A2(_2867_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6404_ (.A1(_0687_),
    .A2(_2956_),
    .B(_3024_),
    .C(_2855_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6405_ (.A1(_1831_),
    .A2(_2856_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6406_ (.A1(\mod.ins_ldr_3 ),
    .A2(_2995_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6407_ (.A1(_3025_),
    .A2(_3026_),
    .B(_3023_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6408_ (.A1(\mod.rd_3[0] ),
    .A2(_2884_),
    .B(_3017_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6409_ (.A1(_1850_),
    .A2(_2883_),
    .B(_3027_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6410_ (.A1(\mod.rd_3[1] ),
    .A2(_2884_),
    .B(_3017_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6411_ (.A1(_1849_),
    .A2(_2883_),
    .B(_3028_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6412_ (.I(_2141_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6413_ (.A1(\mod.rd_3[2] ),
    .A2(_2858_),
    .B(_2140_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6414_ (.A1(_3029_),
    .A2(_2956_),
    .B(_3030_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6415_ (.A1(\mod.rd_3[3] ),
    .A2(_2858_),
    .B(_2140_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6416_ (.A1(_2147_),
    .A2(_2956_),
    .B(_3031_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6417_ (.A1(_2728_),
    .A2(_1801_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6418_ (.I(_3032_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6419_ (.A1(_1812_),
    .A2(_0003_),
    .A3(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6420_ (.I(_3034_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(_1813_),
    .A2(_3033_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6422_ (.I(_1854_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6423_ (.A1(\mod.instr_2[6] ),
    .A2(_3025_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6424_ (.I(_3037_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6425_ (.A1(_3029_),
    .A2(_3036_),
    .A3(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6426_ (.A1(_3035_),
    .A2(_3039_),
    .B(_3023_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6427_ (.A1(_1814_),
    .A2(_3033_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6428_ (.I(_1858_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6429_ (.A1(_3029_),
    .A2(_3041_),
    .A3(_3038_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6430_ (.A1(_3040_),
    .A2(_3042_),
    .B(_3023_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6431_ (.A1(_1815_),
    .A2(_3033_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6432_ (.I(_1852_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6433_ (.A1(_3029_),
    .A2(_3044_),
    .A3(_3038_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6434_ (.I(_2715_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6435_ (.A1(_3043_),
    .A2(_3045_),
    .B(_3046_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6436_ (.I(_3032_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6437_ (.A1(_1825_),
    .A2(_3047_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6438_ (.A1(_2967_),
    .A2(_1862_),
    .A3(_3038_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6439_ (.A1(_3048_),
    .A2(_3049_),
    .B(_3046_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6440_ (.A1(_1824_),
    .A2(_3047_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6441_ (.A1(_2967_),
    .A2(_3036_),
    .A3(_3037_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6442_ (.A1(_3050_),
    .A2(_3051_),
    .B(_3046_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6443_ (.A1(_1822_),
    .A2(_3047_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6444_ (.A1(_2967_),
    .A2(_3041_),
    .A3(_3037_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6445_ (.A1(_3052_),
    .A2(_3053_),
    .B(_3046_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6446_ (.A1(_1826_),
    .A2(_3047_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6447_ (.I(_2966_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6448_ (.A1(_3055_),
    .A2(_3044_),
    .A3(_3037_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6449_ (.I(_2715_),
    .Z(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6450_ (.A1(_3054_),
    .A2(_3056_),
    .B(_3057_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6451_ (.I(_3032_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6452_ (.A1(_2147_),
    .A2(_2966_),
    .A3(_3025_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6453_ (.A1(_1807_),
    .A2(_3058_),
    .B1(_3059_),
    .B2(_1862_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6454_ (.A1(_2992_),
    .A2(_3060_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6455_ (.A1(_1804_),
    .A2(_3058_),
    .B1(_3059_),
    .B2(_3036_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6456_ (.A1(_2992_),
    .A2(_3061_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6457_ (.A1(_1810_),
    .A2(_3058_),
    .B1(_3059_),
    .B2(_3041_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6458_ (.A1(_2716_),
    .A2(_3062_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6459_ (.A1(_1802_),
    .A2(_3058_),
    .B1(_3059_),
    .B2(_3044_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6460_ (.A1(_2716_),
    .A2(_3063_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6461_ (.I(_3032_),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6462_ (.A1(_1817_),
    .A2(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6463_ (.A1(_2147_),
    .A2(_3025_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6464_ (.A1(_3055_),
    .A2(_1862_),
    .A3(_3066_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6465_ (.A1(_3065_),
    .A2(_3067_),
    .B(_3057_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6466_ (.A1(_1818_),
    .A2(_3064_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6467_ (.A1(_3055_),
    .A2(_3036_),
    .A3(_3066_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6468_ (.A1(_3068_),
    .A2(_3069_),
    .B(_3057_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6469_ (.A1(_1819_),
    .A2(_3064_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6470_ (.A1(_3055_),
    .A2(_3041_),
    .A3(_3066_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6471_ (.A1(_3070_),
    .A2(_3071_),
    .B(_3057_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6472_ (.A1(_1820_),
    .A2(_3064_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6473_ (.A1(_2966_),
    .A2(_3044_),
    .A3(_3066_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6474_ (.A1(_3072_),
    .A2(_3073_),
    .B(_2789_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6475_ (.A1(\mod.des.des_counter[0] ),
    .A2(\mod.des.des_counter[1] ),
    .A3(\mod.des.des_counter[2] ),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6476_ (.I(_3074_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6477_ (.I0(\mod.des.des_dout[0] ),
    .I1(net16),
    .S(_3075_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6478_ (.I(_3076_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6479_ (.I0(\mod.des.des_dout[1] ),
    .I1(net17),
    .S(_3075_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6480_ (.I(_3077_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6481_ (.I0(\mod.des.des_dout[2] ),
    .I1(net18),
    .S(_3075_),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6482_ (.I(_3078_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6483_ (.I0(\mod.des.des_dout[3] ),
    .I1(net19),
    .S(_3075_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6484_ (.I(_3079_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6485_ (.I(_3074_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6486_ (.I0(\mod.des.des_dout[4] ),
    .I1(net2),
    .S(_3080_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6487_ (.I(_3081_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6488_ (.I0(\mod.des.des_dout[5] ),
    .I1(net3),
    .S(_3080_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6489_ (.I(_3082_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6490_ (.I0(\mod.des.des_dout[6] ),
    .I1(net4),
    .S(_3080_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6491_ (.I(_3083_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6492_ (.I0(\mod.des.des_dout[7] ),
    .I1(net5),
    .S(_3080_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6493_ (.I(_3084_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6494_ (.I(_3074_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6495_ (.I0(\mod.des.des_dout[8] ),
    .I1(net6),
    .S(_3085_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6496_ (.I(_3086_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6497_ (.I0(\mod.des.des_dout[9] ),
    .I1(net7),
    .S(_3085_),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6498_ (.I(_3087_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6499_ (.I0(\mod.des.des_dout[10] ),
    .I1(net8),
    .S(_3085_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6500_ (.I(_3088_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6501_ (.I0(\mod.des.des_dout[11] ),
    .I1(net9),
    .S(_3085_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6502_ (.I(_3089_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6503_ (.I0(\mod.des.des_dout[12] ),
    .I1(net10),
    .S(_3074_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6504_ (.I(_3090_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6505_ (.A1(_2327_),
    .A2(_2624_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6506_ (.I(_3091_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6507_ (.I(_3092_),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6508_ (.I(_3091_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6509_ (.I(_3094_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6510_ (.A1(\mod.registers.r15[0] ),
    .A2(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6511_ (.A1(_2385_),
    .A2(_3093_),
    .B(_3096_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6512_ (.A1(\mod.registers.r15[1] ),
    .A2(_3095_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6513_ (.A1(_2393_),
    .A2(_3093_),
    .B(_3097_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6514_ (.A1(\mod.registers.r15[2] ),
    .A2(_3095_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6515_ (.A1(_2396_),
    .A2(_3093_),
    .B(_3098_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6516_ (.A1(\mod.registers.r15[3] ),
    .A2(_3095_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6517_ (.A1(_2399_),
    .A2(_3093_),
    .B(_3099_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6518_ (.I(_3092_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6519_ (.I(_3094_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(\mod.registers.r15[4] ),
    .A2(_3101_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6521_ (.A1(_2402_),
    .A2(_3100_),
    .B(_3102_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6522_ (.A1(\mod.registers.r15[5] ),
    .A2(_3101_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6523_ (.A1(_2407_),
    .A2(_3100_),
    .B(_3103_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6524_ (.A1(\mod.registers.r15[6] ),
    .A2(_3101_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6525_ (.A1(_2410_),
    .A2(_3100_),
    .B(_3104_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6526_ (.A1(\mod.registers.r15[7] ),
    .A2(_3101_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6527_ (.A1(_2413_),
    .A2(_3100_),
    .B(_3105_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6528_ (.I(_3092_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6529_ (.I(_3094_),
    .Z(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6530_ (.A1(\mod.registers.r15[8] ),
    .A2(_3107_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6531_ (.A1(_2416_),
    .A2(_3106_),
    .B(_3108_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6532_ (.A1(\mod.registers.r15[9] ),
    .A2(_3107_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6533_ (.A1(_2421_),
    .A2(_3106_),
    .B(_3109_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6534_ (.A1(\mod.registers.r15[10] ),
    .A2(_3107_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6535_ (.A1(_2424_),
    .A2(_3106_),
    .B(_3110_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6536_ (.A1(\mod.registers.r15[11] ),
    .A2(_3107_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6537_ (.A1(_2427_),
    .A2(_3106_),
    .B(_3111_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6538_ (.I(_3092_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6539_ (.I(_3094_),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6540_ (.A1(\mod.registers.r15[12] ),
    .A2(_3113_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6541_ (.A1(_2430_),
    .A2(_3112_),
    .B(_3114_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6542_ (.A1(\mod.registers.r15[13] ),
    .A2(_3113_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6543_ (.A1(_2435_),
    .A2(_3112_),
    .B(_3115_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6544_ (.A1(\mod.registers.r15[14] ),
    .A2(_3113_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6545_ (.A1(_2438_),
    .A2(_3112_),
    .B(_3116_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6546_ (.A1(\mod.registers.r15[15] ),
    .A2(_3113_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6547_ (.A1(_2441_),
    .A2(_3112_),
    .B(_3117_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6548_ (.A1(\mod.des.des_counter[2] ),
    .A2(_1906_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6549_ (.I(_3118_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6550_ (.I0(\mod.des.des_dout[13] ),
    .I1(net16),
    .S(_3119_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6551_ (.I(_3120_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6552_ (.I0(\mod.des.des_dout[14] ),
    .I1(net17),
    .S(_3119_),
    .Z(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6553_ (.I(_3121_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6554_ (.I0(\mod.des.des_dout[15] ),
    .I1(net18),
    .S(_3119_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6555_ (.I(_3122_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6556_ (.I0(\mod.des.des_dout[16] ),
    .I1(net19),
    .S(_3119_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6557_ (.I(_3123_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6558_ (.I(_3118_),
    .Z(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6559_ (.I0(\mod.des.des_dout[17] ),
    .I1(net2),
    .S(_3124_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6560_ (.I(_3125_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6561_ (.I0(\mod.des.des_dout[18] ),
    .I1(net3),
    .S(_3124_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6562_ (.I(_3126_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6563_ (.I0(\mod.des.des_dout[19] ),
    .I1(net4),
    .S(_3124_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6564_ (.I(_3127_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6565_ (.I0(\mod.des.des_dout[20] ),
    .I1(net5),
    .S(_3124_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6566_ (.I(_3128_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6567_ (.I(_3118_),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6568_ (.I0(\mod.des.des_dout[21] ),
    .I1(net6),
    .S(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6569_ (.I(_3130_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6570_ (.I0(\mod.des.des_dout[22] ),
    .I1(net7),
    .S(_3129_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6571_ (.I(_3131_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6572_ (.I0(\mod.des.des_dout[23] ),
    .I1(net8),
    .S(_3129_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6573_ (.I(_3132_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6574_ (.I0(\mod.des.des_dout[24] ),
    .I1(net9),
    .S(_3129_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6575_ (.I(_3133_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6576_ (.I0(\mod.des.des_dout[25] ),
    .I1(net10),
    .S(_3118_),
    .Z(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6577_ (.I(_3134_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6578_ (.A1(\mod.des.des_counter[2] ),
    .A2(_2071_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6579_ (.I(_3135_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6580_ (.I(_3136_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6581_ (.I0(net16),
    .I1(\mod.des.des_dout[26] ),
    .S(_3137_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6582_ (.I(_3138_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6583_ (.I0(net17),
    .I1(\mod.des.des_dout[27] ),
    .S(_3137_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6584_ (.I(_3139_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6585_ (.I0(net18),
    .I1(\mod.des.des_dout[28] ),
    .S(_3137_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6586_ (.I(_3140_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6587_ (.I0(net19),
    .I1(\mod.des.des_dout[29] ),
    .S(_3137_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6588_ (.I(_3141_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6589_ (.I(_3135_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6590_ (.I0(net2),
    .I1(\mod.des.des_dout[30] ),
    .S(_3142_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6591_ (.I(_3143_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6592_ (.I0(net3),
    .I1(\mod.des.des_dout[31] ),
    .S(_3142_),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6593_ (.I(_3144_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6594_ (.I0(net4),
    .I1(\mod.des.des_dout[32] ),
    .S(_3142_),
    .Z(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6595_ (.I(_3145_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6596_ (.I0(net5),
    .I1(\mod.des.des_dout[33] ),
    .S(_3142_),
    .Z(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6597_ (.I(_3146_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6598_ (.I0(net6),
    .I1(\mod.des.des_dout[34] ),
    .S(_3136_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6599_ (.I(_3147_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6600_ (.I0(net7),
    .I1(\mod.des.des_dout[35] ),
    .S(_3136_),
    .Z(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6601_ (.I(_3148_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6602_ (.I0(net8),
    .I1(\mod.des.des_dout[36] ),
    .S(_3136_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6603_ (.I(_3149_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6604_ (.D(_0108_),
    .RN(_0003_),
    .CLK(net218),
    .Q(\mod.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6605_ (.D(_0109_),
    .CLK(net84),
    .Q(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6606_ (.D(_0110_),
    .CLK(net84),
    .Q(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6607_ (.D(_0111_),
    .CLK(net159),
    .Q(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6608_ (.D(_0112_),
    .CLK(net86),
    .Q(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6609_ (.D(_0113_),
    .CLK(net85),
    .Q(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6610_ (.D(_0114_),
    .CLK(net77),
    .Q(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6611_ (.D(_0115_),
    .CLK(net77),
    .Q(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6612_ (.D(_0116_),
    .CLK(net76),
    .Q(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6613_ (.D(_0117_),
    .CLK(net131),
    .Q(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6614_ (.D(_0118_),
    .CLK(net130),
    .Q(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6615_ (.D(_0119_),
    .CLK(net131),
    .Q(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6616_ (.D(_0120_),
    .CLK(net130),
    .Q(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6617_ (.D(_0121_),
    .CLK(net135),
    .Q(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6618_ (.D(_0122_),
    .CLK(net138),
    .Q(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6619_ (.D(_0123_),
    .CLK(net135),
    .Q(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6620_ (.D(_0124_),
    .CLK(net134),
    .Q(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6621_ (.D(_0125_),
    .CLK(net159),
    .Q(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6622_ (.D(_0126_),
    .CLK(net161),
    .Q(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6623_ (.D(_0127_),
    .CLK(net161),
    .Q(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6624_ (.D(_0128_),
    .CLK(net87),
    .Q(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6625_ (.D(_0129_),
    .CLK(net85),
    .Q(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6626_ (.D(_0130_),
    .CLK(net71),
    .Q(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6627_ (.D(_0131_),
    .CLK(net74),
    .Q(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6628_ (.D(_0132_),
    .CLK(net76),
    .Q(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6629_ (.D(_0133_),
    .CLK(net126),
    .Q(\mod.registers.r2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6630_ (.D(_0134_),
    .CLK(net128),
    .Q(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6631_ (.D(_0135_),
    .CLK(net130),
    .Q(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6632_ (.D(_0136_),
    .CLK(net126),
    .Q(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6633_ (.D(_0137_),
    .CLK(net140),
    .Q(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6634_ (.D(_0138_),
    .CLK(net140),
    .Q(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6635_ (.D(_0139_),
    .CLK(net141),
    .Q(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6636_ (.D(_0140_),
    .CLK(net142),
    .Q(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6637_ (.D(_0141_),
    .CLK(net84),
    .Q(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6638_ (.D(_0142_),
    .CLK(net87),
    .Q(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6639_ (.D(_0143_),
    .CLK(net84),
    .Q(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6640_ (.D(_0144_),
    .CLK(net129),
    .Q(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6641_ (.D(_0145_),
    .CLK(net85),
    .Q(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6642_ (.D(_0146_),
    .CLK(net70),
    .Q(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6643_ (.D(_0147_),
    .CLK(net76),
    .Q(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6644_ (.D(_0148_),
    .CLK(net79),
    .Q(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6645_ (.D(_0149_),
    .CLK(net130),
    .Q(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6646_ (.D(_0150_),
    .CLK(net131),
    .Q(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6647_ (.D(_0151_),
    .CLK(net127),
    .Q(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6648_ (.D(_0152_),
    .CLK(net127),
    .Q(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6649_ (.D(_0153_),
    .CLK(net138),
    .Q(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6650_ (.D(_0154_),
    .CLK(net138),
    .Q(\mod.registers.r3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6651_ (.D(_0155_),
    .CLK(net138),
    .Q(\mod.registers.r3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6652_ (.D(_0156_),
    .CLK(net134),
    .Q(\mod.registers.r3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6653_ (.D(_0157_),
    .CLK(net159),
    .Q(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6654_ (.D(_0158_),
    .CLK(net160),
    .Q(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6655_ (.D(_0159_),
    .CLK(net159),
    .Q(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6656_ (.D(_0160_),
    .CLK(net128),
    .Q(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6657_ (.D(_0161_),
    .CLK(net85),
    .Q(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6658_ (.D(_0162_),
    .CLK(net76),
    .Q(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6659_ (.D(_0163_),
    .CLK(net80),
    .Q(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6660_ (.D(_0164_),
    .CLK(net77),
    .Q(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6661_ (.D(_0165_),
    .CLK(net129),
    .Q(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6662_ (.D(_0166_),
    .CLK(net128),
    .Q(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6663_ (.D(_0167_),
    .CLK(net132),
    .Q(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6664_ (.D(_0168_),
    .CLK(net128),
    .Q(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6665_ (.D(_0169_),
    .CLK(net140),
    .Q(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6666_ (.D(_0170_),
    .CLK(net140),
    .Q(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6667_ (.D(_0171_),
    .CLK(net142),
    .Q(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6668_ (.D(_0172_),
    .CLK(net142),
    .Q(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6669_ (.D(_0173_),
    .CLK(net52),
    .Q(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6670_ (.D(_0174_),
    .CLK(net52),
    .Q(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6671_ (.D(_0175_),
    .CLK(net53),
    .Q(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6672_ (.D(_0176_),
    .CLK(net53),
    .Q(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6673_ (.D(_0177_),
    .CLK(net48),
    .Q(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6674_ (.D(_0178_),
    .CLK(net40),
    .Q(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6675_ (.D(_0179_),
    .CLK(net47),
    .Q(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6676_ (.D(_0180_),
    .CLK(net48),
    .Q(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6677_ (.D(_0181_),
    .CLK(net91),
    .Q(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6678_ (.D(_0182_),
    .CLK(net90),
    .Q(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6679_ (.D(_0183_),
    .CLK(net95),
    .Q(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6680_ (.D(_0184_),
    .CLK(net95),
    .Q(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6681_ (.D(_0185_),
    .CLK(net114),
    .Q(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6682_ (.D(_0186_),
    .CLK(net96),
    .Q(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6683_ (.D(_0187_),
    .CLK(net114),
    .Q(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6684_ (.D(_0188_),
    .CLK(net114),
    .Q(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6685_ (.D(_0189_),
    .CLK(net52),
    .Q(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6686_ (.D(_0190_),
    .CLK(net48),
    .Q(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6687_ (.D(_0191_),
    .CLK(net53),
    .Q(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6688_ (.D(_0192_),
    .CLK(net90),
    .Q(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6689_ (.D(_0193_),
    .CLK(net47),
    .Q(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6690_ (.D(_0194_),
    .CLK(net40),
    .Q(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6691_ (.D(_0195_),
    .CLK(net47),
    .Q(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6692_ (.D(_0196_),
    .CLK(net47),
    .Q(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6693_ (.D(_0197_),
    .CLK(net91),
    .Q(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6694_ (.D(_0198_),
    .CLK(net90),
    .Q(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6695_ (.D(_0199_),
    .CLK(net95),
    .Q(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6696_ (.D(_0200_),
    .CLK(net91),
    .Q(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6697_ (.D(_0201_),
    .CLK(net111),
    .Q(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6698_ (.D(_0202_),
    .CLK(net98),
    .Q(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6699_ (.D(_0203_),
    .CLK(net111),
    .Q(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6700_ (.D(_0204_),
    .CLK(net113),
    .Q(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6701_ (.D(_0205_),
    .CLK(net54),
    .Q(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6702_ (.D(_0206_),
    .CLK(net49),
    .Q(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6703_ (.D(_0207_),
    .CLK(net55),
    .Q(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6704_ (.D(_0208_),
    .CLK(net92),
    .Q(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6705_ (.D(_0209_),
    .CLK(net52),
    .Q(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6706_ (.D(_0210_),
    .CLK(net39),
    .Q(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6707_ (.D(_0211_),
    .CLK(net49),
    .Q(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6708_ (.D(_0212_),
    .CLK(net50),
    .Q(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6709_ (.D(_0213_),
    .CLK(net91),
    .Q(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6710_ (.D(_0214_),
    .CLK(net90),
    .Q(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6711_ (.D(_0215_),
    .CLK(net96),
    .Q(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6712_ (.D(_0216_),
    .CLK(net95),
    .Q(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6713_ (.D(_0217_),
    .CLK(net111),
    .Q(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6714_ (.D(_0218_),
    .CLK(net96),
    .Q(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6715_ (.D(_0219_),
    .CLK(net111),
    .Q(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6716_ (.D(_0220_),
    .CLK(net113),
    .Q(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6717_ (.D(_0221_),
    .CLK(net55),
    .Q(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6718_ (.D(_0222_),
    .CLK(net49),
    .Q(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6719_ (.D(_0223_),
    .CLK(net54),
    .Q(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6720_ (.D(_0224_),
    .CLK(net92),
    .Q(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6721_ (.D(_0225_),
    .CLK(net50),
    .Q(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6722_ (.D(_0226_),
    .CLK(net39),
    .Q(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6723_ (.D(_0227_),
    .CLK(net39),
    .Q(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6724_ (.D(_0228_),
    .CLK(net49),
    .Q(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6725_ (.D(_0229_),
    .CLK(net92),
    .Q(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6726_ (.D(_0230_),
    .CLK(net92),
    .Q(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6727_ (.D(_0231_),
    .CLK(net97),
    .Q(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6728_ (.D(_0232_),
    .CLK(net93),
    .Q(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6729_ (.D(_0233_),
    .CLK(net112),
    .Q(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6730_ (.D(_0234_),
    .CLK(net97),
    .Q(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6731_ (.D(_0235_),
    .CLK(net112),
    .Q(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6732_ (.D(_0236_),
    .CLK(net113),
    .Q(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6733_ (.D(_0237_),
    .CLK(net62),
    .Q(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6734_ (.D(_0238_),
    .CLK(net58),
    .Q(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6735_ (.D(_0239_),
    .CLK(net63),
    .Q(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6736_ (.D(_0240_),
    .CLK(net62),
    .Q(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6737_ (.D(_0241_),
    .CLK(net45),
    .Q(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6738_ (.D(_0242_),
    .CLK(net69),
    .Q(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6739_ (.D(_0243_),
    .CLK(net69),
    .Q(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6740_ (.D(_0244_),
    .CLK(net68),
    .Q(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6741_ (.D(_0245_),
    .CLK(net107),
    .Q(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6742_ (.D(_0246_),
    .CLK(net103),
    .Q(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6743_ (.D(_0247_),
    .CLK(net108),
    .Q(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6744_ (.D(_0248_),
    .CLK(net107),
    .Q(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6745_ (.D(_0249_),
    .CLK(net121),
    .Q(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6746_ (.D(_0250_),
    .CLK(net117),
    .Q(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6747_ (.D(_0251_),
    .CLK(net120),
    .Q(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6748_ (.D(_0252_),
    .CLK(net120),
    .Q(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6749_ (.D(_0253_),
    .CLK(net42),
    .Q(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6750_ (.D(_0254_),
    .CLK(net42),
    .Q(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6751_ (.D(_0255_),
    .CLK(net42),
    .Q(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6752_ (.D(_0256_),
    .CLK(net57),
    .Q(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6753_ (.D(_0257_),
    .CLK(net69),
    .Q(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6754_ (.D(_0258_),
    .CLK(net70),
    .Q(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6755_ (.D(_0259_),
    .CLK(net70),
    .Q(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6756_ (.D(_0260_),
    .CLK(net70),
    .Q(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6757_ (.D(_0261_),
    .CLK(net106),
    .Q(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6758_ (.D(_0262_),
    .CLK(net101),
    .Q(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6759_ (.D(_0263_),
    .CLK(net105),
    .Q(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6760_ (.D(_0264_),
    .CLK(net102),
    .Q(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6761_ (.D(_0265_),
    .CLK(net121),
    .Q(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6762_ (.D(_0266_),
    .CLK(net136),
    .Q(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6763_ (.D(_0267_),
    .CLK(net136),
    .Q(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6764_ (.D(_0268_),
    .CLK(net121),
    .Q(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6765_ (.D(_0269_),
    .CLK(net57),
    .Q(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6766_ (.D(_0270_),
    .CLK(net60),
    .Q(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6767_ (.D(_0271_),
    .CLK(net57),
    .Q(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6768_ (.D(_0272_),
    .CLK(net57),
    .Q(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6769_ (.D(_0273_),
    .CLK(net73),
    .Q(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6770_ (.D(_0274_),
    .CLK(net71),
    .Q(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6771_ (.D(_0275_),
    .CLK(net74),
    .Q(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6772_ (.D(_0276_),
    .CLK(net71),
    .Q(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6773_ (.D(_0277_),
    .CLK(net126),
    .Q(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6774_ (.D(_0278_),
    .CLK(net103),
    .Q(\mod.registers.r11[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6775_ (.D(_0279_),
    .CLK(net104),
    .Q(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6776_ (.D(_0280_),
    .CLK(net126),
    .Q(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6777_ (.D(_0281_),
    .CLK(net134),
    .Q(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6778_ (.D(_0282_),
    .CLK(net136),
    .Q(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6779_ (.D(_0283_),
    .CLK(net136),
    .Q(\mod.registers.r11[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6780_ (.D(_0284_),
    .CLK(net134),
    .Q(\mod.registers.r11[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6781_ (.D(_0285_),
    .CLK(net43),
    .Q(\mod.registers.r12[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6782_ (.D(_0286_),
    .CLK(net43),
    .Q(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6783_ (.D(_0287_),
    .CLK(net44),
    .Q(\mod.registers.r12[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6784_ (.D(_0288_),
    .CLK(net43),
    .Q(\mod.registers.r12[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6785_ (.D(_0289_),
    .CLK(net45),
    .Q(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6786_ (.D(_0290_),
    .CLK(net68),
    .Q(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6787_ (.D(_0291_),
    .CLK(net68),
    .Q(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6788_ (.D(_0292_),
    .CLK(net68),
    .Q(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6789_ (.D(_0293_),
    .CLK(net103),
    .Q(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6790_ (.D(_0294_),
    .CLK(net103),
    .Q(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6791_ (.D(_0295_),
    .CLK(net107),
    .Q(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6792_ (.D(_0296_),
    .CLK(net107),
    .Q(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6793_ (.D(_0297_),
    .CLK(net118),
    .Q(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6794_ (.D(_0298_),
    .CLK(net117),
    .Q(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6795_ (.D(_0299_),
    .CLK(net117),
    .Q(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6796_ (.D(_0300_),
    .CLK(net120),
    .Q(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6797_ (.D(_0301_),
    .CLK(net64),
    .Q(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6798_ (.D(_0302_),
    .CLK(net59),
    .Q(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6799_ (.D(_0303_),
    .CLK(net64),
    .Q(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6800_ (.D(_0304_),
    .CLK(net65),
    .Q(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6801_ (.D(_0305_),
    .CLK(net73),
    .Q(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6802_ (.D(_0306_),
    .CLK(net43),
    .Q(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6803_ (.D(_0307_),
    .CLK(net73),
    .Q(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6804_ (.D(_0308_),
    .CLK(net73),
    .Q(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6805_ (.D(_0309_),
    .CLK(net105),
    .Q(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6806_ (.D(_0310_),
    .CLK(net101),
    .Q(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6807_ (.D(_0311_),
    .CLK(net106),
    .Q(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6808_ (.D(_0312_),
    .CLK(net101),
    .Q(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6809_ (.D(_0313_),
    .CLK(net118),
    .Q(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6810_ (.D(_0314_),
    .CLK(net117),
    .Q(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6811_ (.D(_0315_),
    .CLK(net120),
    .Q(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6812_ (.D(_0316_),
    .CLK(net122),
    .Q(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6813_ (.D(_0317_),
    .CLK(net62),
    .Q(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6814_ (.D(_0318_),
    .CLK(net58),
    .Q(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6815_ (.D(_0319_),
    .CLK(net62),
    .Q(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6816_ (.D(_0320_),
    .CLK(net63),
    .Q(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6817_ (.D(_0321_),
    .CLK(net41),
    .Q(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6818_ (.D(_0322_),
    .CLK(net40),
    .Q(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6819_ (.D(_0323_),
    .CLK(net41),
    .Q(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6820_ (.D(_0324_),
    .CLK(net39),
    .Q(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6821_ (.D(_0325_),
    .CLK(net97),
    .Q(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6822_ (.D(_0326_),
    .CLK(net93),
    .Q(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6823_ (.D(_0327_),
    .CLK(net98),
    .Q(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6824_ (.D(_0328_),
    .CLK(net97),
    .Q(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6825_ (.D(_0329_),
    .CLK(net119),
    .Q(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6826_ (.D(_0330_),
    .CLK(net105),
    .Q(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6827_ (.D(_0331_),
    .CLK(net122),
    .Q(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6828_ (.D(_0332_),
    .CLK(net122),
    .Q(\mod.registers.r14[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6829_ (.D(_0000_),
    .SETN(_0004_),
    .CLK(net218),
    .Q(\mod.des.des_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6830_ (.D(_0001_),
    .SETN(_0005_),
    .CLK(net219),
    .Q(\mod.des.des_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _6831_ (.D(_0002_),
    .SETN(_0006_),
    .CLK(net217),
    .Q(\mod.des.des_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6832_ (.D(_0333_),
    .CLK(net176),
    .Q(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6833_ (.D(_0334_),
    .CLK(net175),
    .Q(\mod.valid1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6834_ (.D(_0335_),
    .CLK(net190),
    .Q(\mod.pc0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6835_ (.D(_0336_),
    .CLK(net190),
    .Q(\mod.pc0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6836_ (.D(_0337_),
    .CLK(net180),
    .Q(\mod.pc0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6837_ (.D(_0338_),
    .CLK(net177),
    .Q(\mod.pc0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6838_ (.D(_0339_),
    .CLK(net181),
    .Q(\mod.pc0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6839_ (.D(_0340_),
    .CLK(net177),
    .Q(\mod.pc0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6840_ (.D(_0341_),
    .CLK(net180),
    .Q(\mod.pc0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6841_ (.D(_0342_),
    .CLK(net180),
    .Q(\mod.pc0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6842_ (.D(_0343_),
    .CLK(net186),
    .Q(\mod.pc0[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6843_ (.D(_0344_),
    .CLK(net188),
    .Q(\mod.pc0[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6844_ (.D(_0345_),
    .CLK(net181),
    .Q(\mod.pc0[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6845_ (.D(_0346_),
    .CLK(net189),
    .Q(\mod.pc0[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6846_ (.D(_0347_),
    .CLK(net178),
    .Q(\mod.pc0[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6847_ (.D(_0348_),
    .CLK(net190),
    .Q(\mod.pc0[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6848_ (.D(_0349_),
    .CLK(net198),
    .Q(\mod.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6849_ (.D(_0350_),
    .CLK(net192),
    .Q(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6850_ (.D(_0351_),
    .CLK(net192),
    .Q(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6851_ (.D(_0352_),
    .CLK(net198),
    .Q(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6852_ (.D(_0353_),
    .CLK(net198),
    .Q(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6853_ (.D(_0354_),
    .CLK(net199),
    .Q(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6854_ (.D(_0355_),
    .CLK(net198),
    .Q(\mod.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6855_ (.D(_0356_),
    .CLK(net192),
    .Q(\mod.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6856_ (.D(_0357_),
    .CLK(net192),
    .Q(\mod.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6857_ (.D(_0358_),
    .CLK(net191),
    .Q(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6858_ (.D(_0359_),
    .CLK(net190),
    .Q(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6859_ (.D(_0360_),
    .CLK(net191),
    .Q(\mod.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6860_ (.D(_0361_),
    .CLK(net193),
    .Q(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6861_ (.D(_0362_),
    .CLK(net181),
    .Q(\mod.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6862_ (.D(_0363_),
    .CLK(net196),
    .Q(\mod.pc_1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6863_ (.D(_0364_),
    .CLK(net188),
    .Q(\mod.pc_1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6864_ (.D(_0365_),
    .CLK(net195),
    .Q(\mod.pc_1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6865_ (.D(_0366_),
    .CLK(net197),
    .Q(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6866_ (.D(_0367_),
    .CLK(net196),
    .Q(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6867_ (.D(_0368_),
    .CLK(net196),
    .Q(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6868_ (.D(_0369_),
    .CLK(net196),
    .Q(\mod.pc_1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6869_ (.D(_0370_),
    .CLK(net188),
    .Q(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6870_ (.D(_0371_),
    .CLK(net187),
    .Q(\mod.pc_1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6871_ (.D(_0372_),
    .CLK(net186),
    .Q(\mod.pc_1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6872_ (.D(_0373_),
    .CLK(net187),
    .Q(\mod.pc_1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6873_ (.D(_0374_),
    .CLK(net177),
    .Q(\mod.pc_1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6874_ (.D(_0375_),
    .CLK(net178),
    .Q(\mod.pc_1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6875_ (.D(_0376_),
    .CLK(net180),
    .Q(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6876_ (.D(_0377_),
    .CLK(net155),
    .Q(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6877_ (.D(_0378_),
    .CLK(net156),
    .Q(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6878_ (.D(_0379_),
    .CLK(net153),
    .Q(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6879_ (.D(_0380_),
    .CLK(net151),
    .Q(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6880_ (.D(_0381_),
    .CLK(net151),
    .Q(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6881_ (.D(_0382_),
    .CLK(net151),
    .Q(\mod.instr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6882_ (.D(_0383_),
    .CLK(net151),
    .Q(\mod.instr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6883_ (.D(_0384_),
    .CLK(net155),
    .Q(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6884_ (.D(_0385_),
    .CLK(net163),
    .Q(\mod.instr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6885_ (.D(_0386_),
    .CLK(net163),
    .Q(\mod.instr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6886_ (.D(_0387_),
    .CLK(net170),
    .Q(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6887_ (.D(_0388_),
    .CLK(net171),
    .Q(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6888_ (.D(_0389_),
    .CLK(net171),
    .Q(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6889_ (.D(_0390_),
    .CLK(net171),
    .Q(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6890_ (.D(_0391_),
    .CLK(net170),
    .Q(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6891_ (.D(_0392_),
    .CLK(net172),
    .Q(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6892_ (.D(_0393_),
    .CLK(net172),
    .Q(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6893_ (.D(_0394_),
    .CLK(net172),
    .Q(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6894_ (.D(_0395_),
    .CLK(net172),
    .Q(\mod.instr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6895_ (.D(_0396_),
    .CLK(net170),
    .Q(\mod.instr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6896_ (.D(_0397_),
    .CLK(net170),
    .Q(\mod.instr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6897_ (.D(_0398_),
    .CLK(net177),
    .Q(\mod.valid2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6898_ (.D(_0399_),
    .CLK(net164),
    .Q(\mod.instr_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6899_ (.D(_0400_),
    .CLK(net164),
    .Q(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6900_ (.D(_0401_),
    .CLK(net166),
    .Q(\mod.instr_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6901_ (.D(_0402_),
    .CLK(net155),
    .Q(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6902_ (.D(_0403_),
    .CLK(net155),
    .Q(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6903_ (.D(_0404_),
    .CLK(net154),
    .Q(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6904_ (.D(_0405_),
    .CLK(net152),
    .Q(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6905_ (.D(_0406_),
    .CLK(net162),
    .Q(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6906_ (.D(_0407_),
    .CLK(net161),
    .Q(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6907_ (.D(_0408_),
    .CLK(net160),
    .Q(\mod.funct3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6908_ (.D(_0409_),
    .CLK(net161),
    .Q(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6909_ (.D(_0007_),
    .CLK(net149),
    .Q(\mod.instr_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6910_ (.D(_0008_),
    .CLK(net81),
    .Q(\mod.instr_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6911_ (.D(_0009_),
    .CLK(net81),
    .Q(\mod.instr_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6912_ (.D(_0010_),
    .CLK(net80),
    .Q(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6913_ (.D(_0011_),
    .CLK(net80),
    .Q(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6914_ (.D(_0012_),
    .CLK(net80),
    .Q(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6915_ (.D(_0013_),
    .CLK(net81),
    .Q(\mod.instr_2[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6916_ (.D(_0014_),
    .CLK(net149),
    .Q(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6917_ (.D(_0015_),
    .CLK(net156),
    .Q(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6918_ (.D(_0016_),
    .CLK(net154),
    .Q(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6919_ (.D(_0017_),
    .CLK(net187),
    .Q(\mod.pc_2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6920_ (.D(_0018_),
    .CLK(net202),
    .Q(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6921_ (.D(_0019_),
    .CLK(net202),
    .Q(\mod.pc_2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6922_ (.D(_0020_),
    .CLK(net195),
    .Q(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6923_ (.D(_0021_),
    .CLK(net195),
    .Q(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6924_ (.D(_0022_),
    .CLK(net197),
    .Q(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6925_ (.D(_0023_),
    .CLK(net195),
    .Q(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6926_ (.D(_0024_),
    .CLK(net187),
    .Q(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6927_ (.D(_0025_),
    .CLK(net186),
    .Q(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6928_ (.D(_0026_),
    .CLK(net186),
    .Q(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6929_ (.D(_0027_),
    .CLK(net202),
    .Q(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6930_ (.D(_0028_),
    .CLK(net164),
    .Q(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6931_ (.D(_0029_),
    .CLK(net165),
    .Q(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6932_ (.D(_0030_),
    .CLK(net165),
    .Q(\mod.pc_2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6933_ (.D(_0031_),
    .CLK(net164),
    .Q(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6934_ (.D(_0032_),
    .CLK(net175),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6935_ (.D(_0033_),
    .CLK(net175),
    .Q(\mod.ri_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6936_ (.D(_0034_),
    .CLK(net162),
    .Q(\mod.ins_ldr_3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6937_ (.D(_0035_),
    .CLK(net175),
    .Q(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6938_ (.D(_0036_),
    .CLK(net163),
    .Q(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6939_ (.D(_0037_),
    .CLK(net162),
    .Q(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6940_ (.D(_0038_),
    .CLK(net162),
    .Q(\mod.rd_3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6941_ (.D(_0039_),
    .CLK(net154),
    .Q(\mod.ldr_hzd[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6942_ (.D(_0040_),
    .CLK(net152),
    .Q(\mod.ldr_hzd[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6943_ (.D(_0041_),
    .CLK(net154),
    .Q(\mod.ldr_hzd[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6944_ (.D(_0042_),
    .CLK(net152),
    .Q(\mod.ldr_hzd[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6945_ (.D(_0043_),
    .CLK(net77),
    .Q(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6946_ (.D(_0044_),
    .CLK(net78),
    .Q(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6947_ (.D(_0045_),
    .CLK(net147),
    .Q(\mod.ldr_hzd[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6948_ (.D(_0046_),
    .CLK(net147),
    .Q(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6949_ (.D(_0047_),
    .CLK(net149),
    .Q(\mod.ldr_hzd[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6950_ (.D(_0048_),
    .CLK(net149),
    .Q(\mod.ldr_hzd[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6951_ (.D(_0049_),
    .CLK(net150),
    .Q(\mod.ldr_hzd[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6952_ (.D(_0050_),
    .CLK(net152),
    .Q(\mod.ldr_hzd[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6953_ (.D(_0051_),
    .CLK(net147),
    .Q(\mod.ldr_hzd[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6954_ (.D(_0052_),
    .CLK(net148),
    .Q(\mod.ldr_hzd[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6955_ (.D(_0053_),
    .CLK(net147),
    .Q(\mod.ldr_hzd[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6956_ (.D(_0054_),
    .CLK(net148),
    .Q(\mod.ldr_hzd[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6957_ (.D(_0055_),
    .CLK(net219),
    .Q(\mod.des.des_dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6958_ (.D(_0056_),
    .CLK(net215),
    .Q(\mod.des.des_dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6959_ (.D(_0057_),
    .CLK(net213),
    .Q(\mod.des.des_dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6960_ (.D(_0058_),
    .CLK(net213),
    .Q(\mod.des.des_dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6961_ (.D(_0059_),
    .CLK(net208),
    .Q(\mod.des.des_dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6962_ (.D(_0060_),
    .CLK(net208),
    .Q(\mod.des.des_dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6963_ (.D(_0061_),
    .CLK(net208),
    .Q(\mod.des.des_dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6964_ (.D(_0062_),
    .CLK(net212),
    .Q(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6965_ (.D(_0063_),
    .CLK(net219),
    .Q(\mod.des.des_dout[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6966_ (.D(_0064_),
    .CLK(net217),
    .Q(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6967_ (.D(_0065_),
    .CLK(net219),
    .Q(\mod.des.des_dout[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6968_ (.D(_0066_),
    .CLK(net217),
    .Q(\mod.des.des_dout[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6969_ (.D(_0067_),
    .CLK(net217),
    .Q(\mod.des.des_dout[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6970_ (.D(_0068_),
    .CLK(net59),
    .Q(\mod.registers.r15[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6971_ (.D(_0069_),
    .CLK(net60),
    .Q(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6972_ (.D(_0070_),
    .CLK(net59),
    .Q(\mod.registers.r15[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6973_ (.D(_0071_),
    .CLK(net59),
    .Q(\mod.registers.r15[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6974_ (.D(_0072_),
    .CLK(net45),
    .Q(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6975_ (.D(_0073_),
    .CLK(net41),
    .Q(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6976_ (.D(_0074_),
    .CLK(net41),
    .Q(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6977_ (.D(_0075_),
    .CLK(net45),
    .Q(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6978_ (.D(_0076_),
    .CLK(net102),
    .Q(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6979_ (.D(_0077_),
    .CLK(net101),
    .Q(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6980_ (.D(_0078_),
    .CLK(net106),
    .Q(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6981_ (.D(_0079_),
    .CLK(net105),
    .Q(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6982_ (.D(_0080_),
    .CLK(net116),
    .Q(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6983_ (.D(_0081_),
    .CLK(net116),
    .Q(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6984_ (.D(_0082_),
    .CLK(net116),
    .Q(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6985_ (.D(_0083_),
    .CLK(net116),
    .Q(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6986_ (.D(_0084_),
    .CLK(net216),
    .Q(\mod.des.des_dout[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6987_ (.D(_0085_),
    .CLK(net216),
    .Q(\mod.des.des_dout[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6988_ (.D(_0086_),
    .CLK(net216),
    .Q(\mod.des.des_dout[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6989_ (.D(_0087_),
    .CLK(net221),
    .Q(\mod.des.des_dout[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6990_ (.D(_0088_),
    .CLK(net213),
    .Q(\mod.des.des_dout[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6991_ (.D(_0089_),
    .CLK(net214),
    .Q(\mod.des.des_dout[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6992_ (.D(_0090_),
    .CLK(net214),
    .Q(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6993_ (.D(_0091_),
    .CLK(net213),
    .Q(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6994_ (.D(_0092_),
    .CLK(net211),
    .Q(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6995_ (.D(_0093_),
    .CLK(net211),
    .Q(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6996_ (.D(_0094_),
    .CLK(net210),
    .Q(\mod.des.des_dout[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6997_ (.D(_0095_),
    .CLK(net220),
    .Q(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6998_ (.D(_0096_),
    .CLK(net218),
    .Q(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6999_ (.D(_0097_),
    .CLK(net209),
    .Q(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7000_ (.D(_0098_),
    .CLK(net209),
    .Q(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7001_ (.D(_0099_),
    .CLK(net205),
    .Q(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7002_ (.D(_0100_),
    .CLK(net205),
    .Q(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7003_ (.D(_0101_),
    .CLK(net205),
    .Q(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7004_ (.D(_0102_),
    .CLK(net205),
    .Q(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7005_ (.D(_0103_),
    .CLK(net206),
    .Q(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7006_ (.D(_0104_),
    .CLK(net206),
    .Q(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7007_ (.D(_0105_),
    .CLK(net210),
    .Q(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7008_ (.D(_0106_),
    .CLK(net209),
    .Q(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7009_ (.D(_0107_),
    .CLK(net209),
    .Q(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_286 (.ZN(net286));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_287 (.ZN(net287));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_288 (.ZN(net288));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_289 (.ZN(net289));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_290 (.ZN(net290));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_291 (.ZN(net291));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_292 (.ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_293 (.ZN(net293));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_294 (.ZN(net294));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_295 (.ZN(net295));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_296 (.ZN(net296));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_297 (.ZN(net297));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_298 (.ZN(net298));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_299 (.ZN(net299));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_300 (.ZN(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_301 (.ZN(net301));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_302 (.ZN(net302));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_303 (.ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_304 (.ZN(net304));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_305 (.ZN(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_306 (.ZN(net306));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_328 (.ZN(net328));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_329 (.ZN(net329));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_330 (.ZN(net330));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_331 (.ZN(net331));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_332 (.ZN(net332));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_333 (.ZN(net333));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_334 (.ZN(net334));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_335 (.ZN(net335));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_336 (.ZN(net336));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_337 (.ZN(net337));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_338 (.ZN(net338));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_339 (.ZN(net339));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_340 (.ZN(net340));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_341 (.ZN(net341));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_342 (.ZN(net342));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_343 (.ZN(net343));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_344 (.ZN(net344));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_345 (.ZN(net345));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_346 (.ZN(net346));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_347 (.ZN(net347));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_348 (.ZN(net348));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_349 (.ZN(net349));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_350 (.ZN(net350));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_351 (.ZN(net351));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_352 (.ZN(net352));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_353 (.ZN(net353));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_354 (.ZN(net354));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_355 (.ZN(net355));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_356 (.ZN(net356));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_357 (.ZN(net357));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_358 (.ZN(net358));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_359 (.ZN(net359));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_360 (.ZN(net360));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_361 (.ZN(net361));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_362 (.ZN(net362));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_363 (.ZN(net363));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_364 (.ZN(net364));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_365 (.ZN(net365));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_366 (.ZN(net366));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_367 (.ZN(net367));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_368 (.ZN(net368));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_369 (.ZN(net369));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_370 (.ZN(net370));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_371 (.ZN(net371));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_372 (.ZN(net372));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_373 (.ZN(net373));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_374 (.ZN(net374));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_375 (.ZN(net375));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_376 (.ZN(net376));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_377 (.ZN(net377));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_378 (.ZN(net378));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_379 (.ZN(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input2 (.I(io_in[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input3 (.I(io_in[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input4 (.I(io_in[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input5 (.I(io_in[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input9 (.I(io_in[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input10 (.I(io_in[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(io_in[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(io_in[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(io_in[3]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(io_in[4]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input15 (.I(io_in[5]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(io_in[6]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(io_in[7]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(io_in[8]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input19 (.I(io_in[9]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net46),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net44),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net44),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net46),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net67),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net51),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net51),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout49 (.I(net51),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net51),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout51 (.I(net56),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout52 (.I(net54),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net56),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout56 (.I(net66),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout57 (.I(net61),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net61),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout59 (.I(net61),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net61),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net65),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout62 (.I(net64),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net64),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net89),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout68 (.I(net72),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net72),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout70 (.I(net72),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net75),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout73 (.I(net75),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net83),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout76 (.I(net79),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net79),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout79 (.I(net82),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net82),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net88),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout84 (.I(net86),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout85 (.I(net87),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net146),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout90 (.I(net94),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout91 (.I(net94),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout92 (.I(net94),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net100),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout95 (.I(net99),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net99),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout97 (.I(net99),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net100),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout100 (.I(net110),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout101 (.I(net104),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout102 (.I(net104),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout103 (.I(net104),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net109),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net108),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net108),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net110),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout110 (.I(net125),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net115),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout114 (.I(net115),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout115 (.I(net124),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout116 (.I(net119),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout117 (.I(net119),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net123),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout120 (.I(net123),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout121 (.I(net122),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout122 (.I(net123),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net125),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout125 (.I(net145),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout126 (.I(net133),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net133),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout128 (.I(net132),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout129 (.I(net132),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout130 (.I(net131),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout132 (.I(net133),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout133 (.I(net144),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout134 (.I(net137),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout135 (.I(net137),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout136 (.I(net139),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout137 (.I(net139),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout138 (.I(net143),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout139 (.I(net143),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout142 (.I(net143),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout143 (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net146),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net204),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout147 (.I(net150),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net150),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout149 (.I(net150),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net158),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout151 (.I(net153),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout152 (.I(net157),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout153 (.I(net157),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout154 (.I(net156),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout155 (.I(net156),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout156 (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout157 (.I(net158),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout158 (.I(net169),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout159 (.I(net160),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout160 (.I(net168),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout161 (.I(net168),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout162 (.I(net167),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout163 (.I(net167),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout164 (.I(net166),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout165 (.I(net166),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout166 (.I(net167),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout167 (.I(net168),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout168 (.I(net169),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout169 (.I(net185),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout170 (.I(net173),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout171 (.I(net173),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout172 (.I(net174),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout173 (.I(net174),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout174 (.I(net184),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout175 (.I(net176),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout176 (.I(net179),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout177 (.I(net179),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout178 (.I(net179),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout179 (.I(net183),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout180 (.I(net182),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout181 (.I(net182),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout182 (.I(net183),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout183 (.I(net184),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout184 (.I(net185),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout185 (.I(net203),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout186 (.I(net189),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout187 (.I(net189),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout188 (.I(net189),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout189 (.I(net194),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout190 (.I(net193),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout191 (.I(net193),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout192 (.I(net193),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout193 (.I(net194),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout194 (.I(net201),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout195 (.I(net197),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout196 (.I(net197),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout197 (.I(net200),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout198 (.I(net199),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout199 (.I(net200),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout200 (.I(net201),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout201 (.I(net202),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout202 (.I(net203),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout203 (.I(net204),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout204 (.I(\mod.clk ),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout205 (.I(net207),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout206 (.I(net207),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout207 (.I(net208),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout208 (.I(net212),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout209 (.I(net210),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout210 (.I(net211),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout211 (.I(net212),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout212 (.I(net222),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout213 (.I(net215),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net215),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout215 (.I(net216),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout216 (.I(net221),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout217 (.I(net218),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout218 (.I(net220),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout219 (.I(net221),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout220 (.I(net221),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout221 (.I(net222),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout222 (.I(net1),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__B2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__RN (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__B (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__D (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__D (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__D (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__B1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__I (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__B1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__B1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__B1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__B1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A3 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A3 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A4 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__B1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__C (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__B1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__C1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__B1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__B1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__B1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__B1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__B1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__B1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__B1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__B1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__B1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B1 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__B1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A3 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__I (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__I (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__I (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__B1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__B1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__B1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__B2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__B2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A3 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__I (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__B (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__B (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A3 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__B (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__B (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__B2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__I (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__B (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__B (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__B1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__B1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__B1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__B1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__B1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__I (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__C1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__B1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A4 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A4 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__I (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__B (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A4 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A4 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A3 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__I1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__I (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A4 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A3 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__S (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__B (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__I (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__S (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__S (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__I (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__I (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__B1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__B1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__B1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__B1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__B1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__B1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A4 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__B1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__B1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__I (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__I (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__B1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__B1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__B1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__B1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__I (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__B1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__B1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__B2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__B2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__I (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__B1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__B1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__B1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__B1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__B1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__B1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__B1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__B1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__B1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__B1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__B1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A2 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__I (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A3 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A3 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__I (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__B1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__I (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__B2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__B (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A3 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__B1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__B1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__B1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__C (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A3 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__B (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__B (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__B (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__I (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__I (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__B1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__B2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A3 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__B (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__S (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__B (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__C1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__B1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__B1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__C2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__C1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__C1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__C2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__I (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__B1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__I (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__B1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__B1 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__B2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__B2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__C (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A3 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A3 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__B (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__I1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__I1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__C (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__B (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__C (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__B1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__B2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__B (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__I0 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A4 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A4 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__B (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__I0 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A4 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__C (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__B2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A3 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__B (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__I0 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__B1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__B2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__C (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__B2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I0 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__B (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__I1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__B1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__C (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__C (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__B1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__B2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__B (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A3 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A3 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A3 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__B1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__C2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__C1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__B1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__B1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__B1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__B1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__C2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__B1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__B1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__B1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__B1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__B1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__C1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__B1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__C (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__A3 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A3 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__C (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__I1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__B (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__B (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__I (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__B (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__C (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A3 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__B1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A2 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__B1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__B1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__B1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__B1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__C1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__C1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__B1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A3 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A3 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__B1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__B1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__B1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__B1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__B1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__B1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__B1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__B1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__B1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__B1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__B2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__B1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__B1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__B1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__C2 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__B1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__B2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__I (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__B (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__I (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A3 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A3 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A3 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A3 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A3 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A4 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A3 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__B (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__B (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__I (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__B (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__B (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__C (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A4 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__B1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__B2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__I (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__B (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__B (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A3 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A4 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__B1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__B2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A3 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__B (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__C (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__B2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__B1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__B2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__I (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A3 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__B (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A4 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__B (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A3 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A3 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__B (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A3 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A3 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A3 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__B1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__B1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__B1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__B1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__B1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__B1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__B1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__B1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__B1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__C2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__C2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A3 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A3 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__I1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A3 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A4 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A3 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__C (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A3 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__B (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__I (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__B2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__B (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__B (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__B (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__B1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__C (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__I (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__B (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__C (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__B (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__B (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__B2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__C (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__I (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__C (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__C (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__C (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__B1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__C1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__C1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__B1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__B1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__B1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__B1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__B1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__C2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__C1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__B1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__B1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__C1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__B1 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__B1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__C1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__B1 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__B (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__I (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__B (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__B1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__B (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__I (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A4 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A4 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A4 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A4 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A4 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__B (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A3 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A4 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A3 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A3 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A3 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__B1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__B2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__B (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__I (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__I (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A3 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__B1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__C (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__I (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A2 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__I (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A3 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__B1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__B2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A3 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__B (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__I (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A3 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__C (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__B (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__B (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__B (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__I0 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A3 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__B1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__B1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__B (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A3 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A3 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__I (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A3 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__B (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A3 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A3 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A3 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A3 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__B2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A3 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A3 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__B (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__I (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__B (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A3 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A3 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__I (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A3 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__B (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A4 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__B2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__C (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__I (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__C (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__B (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__I (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__B (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__B (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__C (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__B (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__C (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A3 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__B (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__C (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__B (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A1 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__C (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__B (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__B (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__B (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__C (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__B2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__B (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A3 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A3 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__B (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__B (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__B (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__B2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__B2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I0 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I0 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__S (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__S (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__S (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__B2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__B (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I0 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__B (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__C (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__B2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__B2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__B2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__B2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__B (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__B2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__B (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__B2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__B (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__C2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__B (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__B (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__B (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__B (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__B (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__S (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__I0 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__B1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A3 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A3 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__B1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__I (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__C (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__B2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__B1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__B1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__B1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__B2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A3 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A3 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__B (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__I (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__B (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__B (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__C (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__I (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__B3 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__B (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__C (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__B (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I0 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I0 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__B (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__B (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__S (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__I1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I0 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__C (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__B2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__B1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__B (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__C (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__I (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__B (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__B (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__B (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__B (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A3 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A3 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__C (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__B2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A3 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A3 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__B1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__B2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__B2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__B (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__B2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__B (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__B (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__C (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__B (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__B (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__B (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I0 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__S (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__C (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__C (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A3 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A3 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__B1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__B (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__C (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__B1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A3 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A3 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__B1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__B1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__B2 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A4 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A3 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__B1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__B1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B1 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A4 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__B2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__B2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__C1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__B1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__C (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__B (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A3 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__B (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__B1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A4 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A3 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__B (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__C (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__B1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__B1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__B (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__C (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A3 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A3 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__C (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A4 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A4 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__I (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__B (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__B (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__B1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A3 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__C2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__S0 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__S0 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A4 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B2 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__S1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__S1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__B2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__C2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A4 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__C1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I0 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A3 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I3 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__B2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I0 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A3 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__C2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__B2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I3 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__B2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A3 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A4 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__C1 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__B2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__C2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__C2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__C2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__I (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__I (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__B1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__B1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__B1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__C2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__I (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__B1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__B1 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__B2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__I (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A3 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A2 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__S (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__S (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__B (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__C (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__I (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A2 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__I (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__B2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__B2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__B2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__B2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A3 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__C (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__B2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__B1 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__B (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__B (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__B (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__C (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A1 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A3 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__B2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A3 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__B1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__B2 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__B1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__B2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A1 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A3 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__B (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__B (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__C (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A3 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__B1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__B2 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__B1 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__I (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A3 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__B2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A3 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__B1 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__B (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__B2 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A3 (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__I1 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__B1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__C (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__B (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__C (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__B2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__B2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__B2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A1 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__B1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__C (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__B1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__B (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__I (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__C (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__I (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__B (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__I (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__I (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A3 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__I (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A3 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__I (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A3 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__I (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__B (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__B (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__I (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__I (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__B (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__B (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__B (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__I (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__B (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A2 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__B (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__I (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__B1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__B (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__B (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__B (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__I (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__B (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__C (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__B (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__I (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__I (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__B (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__I (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__B1 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__I (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__I (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A1 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__I (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__I (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__I (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__I (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__I (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__I (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__I (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__I (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__I (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__I (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__I (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__I (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A1 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__I (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__I (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__I (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__I (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A2 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A2 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__I (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__I (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__I (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A2 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__I (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__I (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__I (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__I (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__I (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__I (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__I (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__I (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__I (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__I (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__I (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A2 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A2 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A2 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__I (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__I (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__I (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__I (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__I (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A2 (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__I (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__I (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__I (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A2 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A3 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A2 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__I (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__I (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__I (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__I (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__B (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__B (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__I (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__I (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__I (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A3 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__I (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A2 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__I (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__C (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__C (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__C (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__I (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__I (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__I (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__I (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__B (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__B (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__B (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__B (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__I (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__I (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__I (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__I (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__I (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__I (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__I (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__I (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__C (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__C (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__B (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__B (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__B (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__B (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__B (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__B (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__C (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__C (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__C (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__I (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__I (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__B (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__I (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__B (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__B (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__B (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__B (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__B (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__B (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__B (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A2 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A4 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__I (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__I (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__I (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__I (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__I (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__B (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__B (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__B (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__B (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A2 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__I (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__I (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__I (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__B2 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__I (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__I (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__I (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__B2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__B2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__B2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__C (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__C (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__C (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__C (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__B2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__B2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__B2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__B2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__C (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__C (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__C (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__C (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__B2 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__B2 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__B2 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__B2 (.I(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A2 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__C (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__C (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__C (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__C (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__B2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__B2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__B2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__B2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__B2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__B2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__B2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__B2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__B1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__I (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__I (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__I (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__I (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__B1 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__B1 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__B1 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__I (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__I (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__I (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A2 (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__B1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__B1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__B1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A1 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__B (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__B (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__B (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__B (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__B (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__B (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__B (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__B (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__B (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__B (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A3 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__I (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__I (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__I (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__I (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__B2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A3 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A3 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A3 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A3 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__B2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__B (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__B (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__B (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__B (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__B (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__B (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__B (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__B (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__S (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__I (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__I (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__I (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__S (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__S (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__S (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__S (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__S (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__S (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__S (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__S (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__S (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__S (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__S (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__S (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__I (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__I (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__I (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__I (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__I (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__I (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__S (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__I (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__I (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__I (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__S (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__S (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__S (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__S (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__S (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__S (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__S (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__S (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__S (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__S (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__S (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__S (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__I (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__I (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__S (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__S (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__S (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__I (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__S (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__S (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__S (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__S (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__B2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__B2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__B2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A3 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A3 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__I (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__I (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__I (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__B1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__B1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__I (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__I (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__C2 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__B1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A3 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A3 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__I (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__B1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A3 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A3 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__B1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__I (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__B1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__B1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A2 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__I (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A3 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A4 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A4 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A4 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__B1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__B1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__B1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A4 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A4 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__I (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__I (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__I (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__C1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__B1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__B1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__C2 (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__I (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__I (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__C2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__C2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__I (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__B1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__B1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__I (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__I (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__B1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__B1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A2 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__I (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__I (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__B1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__B1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__B1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__B1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__C1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__I (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__I (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__I (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__B1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__I (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__B1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__B1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__I (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__I (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A3 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__B1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__B1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__I (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__B1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__I (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__B1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__B1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__B1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__C (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A3 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A3 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__I0 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__I (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__I (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__I (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A1 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A1 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A2 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__I (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__I (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__B (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__I (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__I (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__I (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__B (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__B (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__I (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__B (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__B (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__I (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__B (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__C (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A3 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A3 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A3 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__C (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__I1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__B (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__I (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__S (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__S (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__I (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__I (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__I (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__C (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A1 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__B (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__B (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__I (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__B (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__I (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__I (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__B (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__I (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__I (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__I (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__B1 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__I (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__B1 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A1 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A3 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__B1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__I (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__I (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__B1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__B1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__A3 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A3 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B1 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__I (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__I (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__B1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__B1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__B1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__I (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__B1 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__I (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__B1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__I0 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(\mod.des.des_dout[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__I0 (.I(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(\mod.des.des_dout[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__I0 (.I(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(\mod.des.des_dout[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__I0 (.I(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(\mod.des.des_dout[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__I0 (.I(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(\mod.des.des_dout[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__I0 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(\mod.des.des_dout[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__I1 (.I(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A1 (.I(\mod.des.des_dout[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__I1 (.I(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(\mod.des.des_dout[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__I1 (.I(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(\mod.des.des_dout[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__I1 (.I(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(\mod.des.des_dout[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__I1 (.I(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(\mod.des.des_dout[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__I1 (.I(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(\mod.des.des_dout[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I1 (.I(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(\mod.des.des_dout[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I1 (.I(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(\mod.des.des_dout[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I1 (.I(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(\mod.des.des_dout[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__I1 (.I(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(\mod.des.des_dout[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__I1 (.I(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A1 (.I(\mod.des.des_dout[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I0 (.I(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(\mod.des.des_dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__I0 (.I(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(\mod.des.des_dout[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A3 (.I(\mod.funct3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__I (.I(\mod.funct3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I1 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I0 (.I(\mod.funct7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__I (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I0 (.I(\mod.funct7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__I (.I(\mod.funct7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__B2 (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__I (.I(\mod.instr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__B2 (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__I (.I(\mod.instr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__B2 (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__I (.I(\mod.instr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__B2 (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(\mod.instr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__B2 (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__I (.I(\mod.instr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__B2 (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__I (.I(\mod.instr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__B2 (.I(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(\mod.instr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__B2 (.I(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I (.I(\mod.instr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__B2 (.I(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__I (.I(\mod.instr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B2 (.I(\mod.instr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__I (.I(\mod.instr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__B2 (.I(\mod.instr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__I (.I(\mod.instr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__B2 (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__I (.I(\mod.instr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B2 (.I(\mod.instr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__I (.I(\mod.instr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__B2 (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I (.I(\mod.instr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B2 (.I(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__I (.I(\mod.instr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__B2 (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__I (.I(\mod.instr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__B2 (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__I (.I(\mod.instr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__I (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A2 (.I(\mod.instr_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__I (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__I (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__I (.I(\mod.instr_2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__I (.I(\mod.instr_2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A2 (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__I (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__I (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__I (.I(\mod.instr_2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__B (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__I (.I(\mod.instr_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__I (.I(\mod.instr_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A1 (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__I (.I(\mod.instr_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__C (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__C (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__I0 (.I(\mod.instr_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(\mod.instr_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(\mod.ldr_hzd[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__B2 (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I (.I(\mod.ldr_hzd[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__C2 (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(\mod.ldr_hzd[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__B (.I(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__I (.I(\mod.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__I (.I(\mod.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__I (.I(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A1 (.I(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(\mod.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__B (.I(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(\mod.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__B (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I (.I(\mod.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__B (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(\mod.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__B (.I(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(\mod.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I0 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(\mod.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(\mod.pc_1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(\mod.pc_1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(\mod.pc_1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(\mod.pc_1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(\mod.pc_1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__I (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(\mod.pc_2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A1 (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A1 (.I(\mod.pc_2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A1 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__I (.I(\mod.pc_2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__I (.I(\mod.pc_2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(\mod.pc_2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(\mod.pc_2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__I (.I(\mod.pc_2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(\mod.pc_2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__I (.I(\mod.pc_2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A1 (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__I (.I(\mod.pc_2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__I (.I(\mod.pc_2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(\mod.rd_3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A1 (.I(\mod.rd_3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(\mod.rd_3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__B2 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(\mod.registers.r10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__B2 (.I(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__B2 (.I(\mod.registers.r10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__B2 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__B2 (.I(\mod.registers.r10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__B2 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__B2 (.I(\mod.registers.r10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__B2 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__B2 (.I(\mod.registers.r10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__C2 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__B2 (.I(\mod.registers.r10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__B2 (.I(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__B2 (.I(\mod.registers.r10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__B2 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__B2 (.I(\mod.registers.r10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__B2 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(\mod.registers.r10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A1 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__B2 (.I(\mod.registers.r10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__C1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A1 (.I(\mod.registers.r10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__B2 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__B2 (.I(\mod.registers.r10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__B2 (.I(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__B2 (.I(\mod.registers.r10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__B2 (.I(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__B2 (.I(\mod.registers.r10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__B2 (.I(\mod.registers.r10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__B2 (.I(\mod.registers.r10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__A1 (.I(\mod.registers.r11[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__B2 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(\mod.registers.r11[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(\mod.registers.r11[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A1 (.I(\mod.registers.r11[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(\mod.registers.r11[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__B2 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A1 (.I(\mod.registers.r11[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A3 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(\mod.registers.r11[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(\mod.registers.r11[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__B2 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__B2 (.I(\mod.registers.r11[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__C2 (.I(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(\mod.registers.r11[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A1 (.I(\mod.registers.r11[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A1 (.I(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(\mod.registers.r11[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__C1 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A3 (.I(\mod.registers.r11[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(\mod.registers.r11[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A3 (.I(\mod.registers.r11[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A1 (.I(\mod.registers.r11[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(\mod.registers.r12[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__B2 (.I(\mod.registers.r12[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__I (.I(\mod.registers.r12[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__B2 (.I(\mod.registers.r12[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__B2 (.I(\mod.registers.r12[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(\mod.registers.r12[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A1 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__B2 (.I(\mod.registers.r12[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__C1 (.I(\mod.registers.r12[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__B2 (.I(\mod.registers.r12[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__B2 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A1 (.I(\mod.registers.r12[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A1 (.I(\mod.registers.r12[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__B2 (.I(\mod.registers.r12[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__B2 (.I(\mod.registers.r12[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__B2 (.I(\mod.registers.r12[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(\mod.registers.r12[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__B2 (.I(\mod.registers.r12[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__A1 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__B2 (.I(\mod.registers.r13[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__B2 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(\mod.registers.r13[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__B2 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A1 (.I(\mod.registers.r13[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__B2 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A1 (.I(\mod.registers.r13[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__B2 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(\mod.registers.r13[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__B2 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(\mod.registers.r13[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A1 (.I(\mod.registers.r13[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A3 (.I(\mod.registers.r13[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A1 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__B2 (.I(\mod.registers.r13[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__B2 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(\mod.registers.r13[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__B2 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A1 (.I(\mod.registers.r13[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__B2 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(\mod.registers.r13[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__B2 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A1 (.I(\mod.registers.r13[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__B2 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(\mod.registers.r13[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__B2 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(\mod.registers.r13[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A3 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(\mod.registers.r13[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__A1 (.I(\mod.registers.r14[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A1 (.I(\mod.registers.r14[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(\mod.registers.r14[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(\mod.registers.r14[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(\mod.registers.r14[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A1 (.I(\mod.registers.r14[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(\mod.registers.r14[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A1 (.I(\mod.registers.r14[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B2 (.I(\mod.registers.r14[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A3 (.I(\mod.registers.r14[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(\mod.registers.r14[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A1 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(\mod.registers.r14[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(\mod.registers.r14[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__B2 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(\mod.registers.r14[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(\mod.registers.r14[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__A1 (.I(\mod.registers.r14[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(\mod.registers.r14[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A3 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(\mod.registers.r14[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(\mod.registers.r15[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A1 (.I(\mod.registers.r15[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__I (.I(\mod.registers.r15[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A1 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A1 (.I(\mod.registers.r15[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(\mod.registers.r15[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__C2 (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__I (.I(\mod.registers.r15[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(\mod.registers.r15[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(\mod.registers.r15[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__B2 (.I(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__B2 (.I(\mod.registers.r15[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__A1 (.I(\mod.registers.r15[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A1 (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__I (.I(\mod.registers.r15[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(\mod.registers.r15[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(\mod.registers.r15[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(\mod.registers.r15[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__B2 (.I(\mod.registers.r15[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A1 (.I(\mod.registers.r15[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__B2 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__B2 (.I(\mod.registers.r1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__B2 (.I(\mod.registers.r1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__B2 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__B2 (.I(\mod.registers.r1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__B2 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__B2 (.I(\mod.registers.r1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__B2 (.I(\mod.registers.r1[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__B2 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__B2 (.I(\mod.registers.r1[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__B2 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A1 (.I(\mod.registers.r1[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__B2 (.I(\mod.registers.r1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__B2 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__B2 (.I(\mod.registers.r1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__B2 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__B2 (.I(\mod.registers.r1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__B2 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__B2 (.I(\mod.registers.r1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__B2 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__B2 (.I(\mod.registers.r1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__B2 (.I(\mod.registers.r1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A3 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__B2 (.I(\mod.registers.r1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A3 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(\mod.registers.r1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__B2 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B2 (.I(\mod.registers.r1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__B2 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__C1 (.I(\mod.registers.r2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__C1 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__B2 (.I(\mod.registers.r2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__C1 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__B2 (.I(\mod.registers.r2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__B2 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B2 (.I(\mod.registers.r2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A1 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__C2 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B2 (.I(\mod.registers.r2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__B2 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__B2 (.I(\mod.registers.r2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__B2 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__C2 (.I(\mod.registers.r2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__B2 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A1 (.I(\mod.registers.r2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A3 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__C1 (.I(\mod.registers.r2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__C1 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__B2 (.I(\mod.registers.r2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A1 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__B2 (.I(\mod.registers.r2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__B2 (.I(\mod.registers.r2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__C1 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__B2 (.I(\mod.registers.r2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__B2 (.I(\mod.registers.r2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__B2 (.I(\mod.registers.r2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__B2 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A1 (.I(\mod.registers.r3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__C1 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__B2 (.I(\mod.registers.r3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__B2 (.I(\mod.registers.r3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__B2 (.I(\mod.registers.r3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__B2 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A1 (.I(\mod.registers.r3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B2 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(\mod.registers.r3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A1 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__B2 (.I(\mod.registers.r3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__B2 (.I(\mod.registers.r3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A1 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__B2 (.I(\mod.registers.r3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__B2 (.I(\mod.registers.r3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__B2 (.I(\mod.registers.r3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__B2 (.I(\mod.registers.r3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__B2 (.I(\mod.registers.r3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A1 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A1 (.I(\mod.registers.r4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__B2 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(\mod.registers.r4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__C2 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A1 (.I(\mod.registers.r4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A1 (.I(\mod.registers.r4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__C1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A1 (.I(\mod.registers.r4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__B2 (.I(\mod.registers.r4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__B2 (.I(\mod.registers.r4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A1 (.I(\mod.registers.r4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A1 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A3 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A1 (.I(\mod.registers.r4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(\mod.registers.r4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__B2 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(\mod.registers.r4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A1 (.I(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(\mod.registers.r4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B2 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(\mod.registers.r4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A3 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A1 (.I(\mod.registers.r4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__B2 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(\mod.registers.r4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A3 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(\mod.registers.r4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__B2 (.I(\mod.registers.r5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(\mod.registers.r5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__B2 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(\mod.registers.r5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__B2 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(\mod.registers.r5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__B2 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(\mod.registers.r5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__B2 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(\mod.registers.r5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__B2 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(\mod.registers.r5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__B2 (.I(\mod.registers.r5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A1 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__B2 (.I(\mod.registers.r5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__B2 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(\mod.registers.r5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(\mod.registers.r5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(\mod.registers.r5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A1 (.I(\mod.registers.r5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__C2 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(\mod.registers.r5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__B2 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(\mod.registers.r5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__B2 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A1 (.I(\mod.registers.r5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__B2 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A1 (.I(\mod.registers.r6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A1 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__B2 (.I(\mod.registers.r6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B2 (.I(\mod.registers.r6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__B2 (.I(\mod.registers.r6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B2 (.I(\mod.registers.r6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__C2 (.I(\mod.registers.r6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A1 (.I(\mod.registers.r6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A1 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__B2 (.I(\mod.registers.r6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B2 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(\mod.registers.r6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__B2 (.I(\mod.registers.r6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__B2 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__B2 (.I(\mod.registers.r6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__B2 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__B2 (.I(\mod.registers.r6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__B2 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__B2 (.I(\mod.registers.r6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__B2 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__B2 (.I(\mod.registers.r6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A1 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__B2 (.I(\mod.registers.r6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__B2 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__B2 (.I(\mod.registers.r6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__B2 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__B2 (.I(\mod.registers.r7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__B2 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__B2 (.I(\mod.registers.r7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__B2 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__B2 (.I(\mod.registers.r7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__B2 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(\mod.registers.r7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__C2 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__B2 (.I(\mod.registers.r7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__B2 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(\mod.registers.r7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__B2 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__B2 (.I(\mod.registers.r7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__B2 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__C1 (.I(\mod.registers.r7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B2 (.I(\mod.registers.r7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__B2 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A1 (.I(\mod.registers.r7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(\mod.registers.r7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__B2 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B2 (.I(\mod.registers.r7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__B2 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__B2 (.I(\mod.registers.r7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A1 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__B2 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__B2 (.I(\mod.registers.r7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__B2 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A1 (.I(\mod.registers.r7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__C2 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__B2 (.I(\mod.registers.r7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__B2 (.I(\mod.registers.r8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__C2 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(\mod.registers.r8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A1 (.I(\mod.registers.r8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__A1 (.I(\mod.registers.r8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__B2 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A1 (.I(\mod.registers.r8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__B2 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__B2 (.I(\mod.registers.r8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__C2 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A1 (.I(\mod.registers.r8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__B2 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A1 (.I(\mod.registers.r8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__B2 (.I(\mod.registers.r8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__B2 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A1 (.I(\mod.registers.r8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__B2 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__B2 (.I(\mod.registers.r8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(\mod.registers.r8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__B2 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(\mod.registers.r8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A3 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(\mod.registers.r8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A3 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A3 (.I(\mod.registers.r8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__C2 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A1 (.I(\mod.registers.r8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__B2 (.I(\mod.registers.r9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__B2 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(\mod.registers.r9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__B2 (.I(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A1 (.I(\mod.registers.r9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__B2 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(\mod.registers.r9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__B2 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(\mod.registers.r9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__C2 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__B2 (.I(\mod.registers.r9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B2 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A1 (.I(\mod.registers.r9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__B2 (.I(\mod.registers.r9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__B2 (.I(\mod.registers.r9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__B2 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(\mod.registers.r9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__C2 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__B2 (.I(\mod.registers.r9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B2 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(\mod.registers.r9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__B2 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(\mod.registers.r9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__B2 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A1 (.I(\mod.registers.r9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__C2 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B2 (.I(\mod.registers.r9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__B2 (.I(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(\mod.registers.r9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__B (.I(\mod.valid0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(\mod.valid_out3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__I1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__I1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__I1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__I0 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__CLK (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__CLK (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__CLK (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__CLK (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__CLK (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__CLK (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__CLK (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__CLK (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__CLK (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__CLK (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__CLK (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__CLK (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__CLK (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__CLK (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__CLK (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__CLK (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__CLK (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__CLK (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__CLK (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__CLK (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__CLK (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout155_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__CLK (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout159_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__CLK (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout166_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout163_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout167_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout160_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout161_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout168_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout158_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout170_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout171_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout172_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout173_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__CLK (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A1 (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout175_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__CLK (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout177_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout178_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout176_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__CLK (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout180_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout181_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout183_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout174_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout184_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout169_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__CLK (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__CLK (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__CLK (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__CLK (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout187_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout188_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout186_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__CLK (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__CLK (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout190_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout191_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout193_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout189_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__CLK (.I(net195));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__CLK (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__CLK (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout200_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout201_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__CLK (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout185_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout203_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__CLK (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout209_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__CLK (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout213_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout214_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__CLK (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout217_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout219_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout220_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout216_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout221_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1044 ();
 assign io_oeb[0] = net223;
 assign io_oeb[10] = net233;
 assign io_oeb[11] = net234;
 assign io_oeb[12] = net235;
 assign io_oeb[13] = net236;
 assign io_oeb[14] = net237;
 assign io_oeb[15] = net238;
 assign io_oeb[16] = net239;
 assign io_oeb[17] = net240;
 assign io_oeb[18] = net241;
 assign io_oeb[19] = net242;
 assign io_oeb[1] = net224;
 assign io_oeb[20] = net243;
 assign io_oeb[21] = net244;
 assign io_oeb[22] = net245;
 assign io_oeb[23] = net246;
 assign io_oeb[24] = net247;
 assign io_oeb[25] = net248;
 assign io_oeb[26] = net249;
 assign io_oeb[27] = net250;
 assign io_oeb[28] = net251;
 assign io_oeb[29] = net252;
 assign io_oeb[2] = net225;
 assign io_oeb[30] = net253;
 assign io_oeb[31] = net254;
 assign io_oeb[32] = net255;
 assign io_oeb[33] = net256;
 assign io_oeb[34] = net257;
 assign io_oeb[35] = net258;
 assign io_oeb[36] = net259;
 assign io_oeb[37] = net260;
 assign io_oeb[3] = net226;
 assign io_oeb[4] = net227;
 assign io_oeb[5] = net228;
 assign io_oeb[6] = net229;
 assign io_oeb[7] = net230;
 assign io_oeb[8] = net231;
 assign io_oeb[9] = net232;
 assign io_out[19] = net261;
 assign io_out[20] = net262;
 assign io_out[21] = net263;
 assign io_out[22] = net264;
 assign io_out[23] = net265;
 assign io_out[24] = net266;
 assign io_out[25] = net267;
 assign io_out[26] = net268;
 assign io_out[27] = net269;
 assign io_out[28] = net270;
 assign io_out[29] = net271;
 assign io_out[30] = net272;
 assign io_out[31] = net273;
 assign io_out[32] = net274;
 assign io_out[33] = net275;
 assign io_out[34] = net276;
 assign io_out[35] = net277;
 assign io_out[36] = net278;
 assign io_out[37] = net279;
 assign la_data_out[0] = net280;
 assign la_data_out[10] = net290;
 assign la_data_out[11] = net291;
 assign la_data_out[12] = net292;
 assign la_data_out[13] = net293;
 assign la_data_out[14] = net294;
 assign la_data_out[15] = net295;
 assign la_data_out[16] = net296;
 assign la_data_out[17] = net297;
 assign la_data_out[18] = net298;
 assign la_data_out[19] = net299;
 assign la_data_out[1] = net281;
 assign la_data_out[20] = net300;
 assign la_data_out[21] = net301;
 assign la_data_out[22] = net302;
 assign la_data_out[23] = net303;
 assign la_data_out[24] = net304;
 assign la_data_out[25] = net305;
 assign la_data_out[26] = net306;
 assign la_data_out[27] = net307;
 assign la_data_out[28] = net308;
 assign la_data_out[29] = net309;
 assign la_data_out[2] = net282;
 assign la_data_out[30] = net310;
 assign la_data_out[31] = net311;
 assign la_data_out[32] = net312;
 assign la_data_out[33] = net313;
 assign la_data_out[34] = net314;
 assign la_data_out[35] = net315;
 assign la_data_out[36] = net316;
 assign la_data_out[37] = net317;
 assign la_data_out[38] = net318;
 assign la_data_out[39] = net319;
 assign la_data_out[3] = net283;
 assign la_data_out[40] = net320;
 assign la_data_out[41] = net321;
 assign la_data_out[42] = net322;
 assign la_data_out[43] = net323;
 assign la_data_out[44] = net324;
 assign la_data_out[45] = net325;
 assign la_data_out[46] = net326;
 assign la_data_out[47] = net327;
 assign la_data_out[48] = net328;
 assign la_data_out[49] = net329;
 assign la_data_out[4] = net284;
 assign la_data_out[50] = net330;
 assign la_data_out[51] = net331;
 assign la_data_out[52] = net332;
 assign la_data_out[53] = net333;
 assign la_data_out[54] = net334;
 assign la_data_out[55] = net335;
 assign la_data_out[56] = net336;
 assign la_data_out[57] = net337;
 assign la_data_out[58] = net338;
 assign la_data_out[59] = net339;
 assign la_data_out[5] = net285;
 assign la_data_out[60] = net340;
 assign la_data_out[61] = net341;
 assign la_data_out[62] = net342;
 assign la_data_out[63] = net343;
 assign la_data_out[6] = net286;
 assign la_data_out[7] = net287;
 assign la_data_out[8] = net288;
 assign la_data_out[9] = net289;
 assign user_irq[0] = net344;
 assign user_irq[1] = net345;
 assign user_irq[2] = net346;
 assign wbs_ack_o = net347;
 assign wbs_dat_o[0] = net348;
 assign wbs_dat_o[10] = net358;
 assign wbs_dat_o[11] = net359;
 assign wbs_dat_o[12] = net360;
 assign wbs_dat_o[13] = net361;
 assign wbs_dat_o[14] = net362;
 assign wbs_dat_o[15] = net363;
 assign wbs_dat_o[16] = net364;
 assign wbs_dat_o[17] = net365;
 assign wbs_dat_o[18] = net366;
 assign wbs_dat_o[19] = net367;
 assign wbs_dat_o[1] = net349;
 assign wbs_dat_o[20] = net368;
 assign wbs_dat_o[21] = net369;
 assign wbs_dat_o[22] = net370;
 assign wbs_dat_o[23] = net371;
 assign wbs_dat_o[24] = net372;
 assign wbs_dat_o[25] = net373;
 assign wbs_dat_o[26] = net374;
 assign wbs_dat_o[27] = net375;
 assign wbs_dat_o[28] = net376;
 assign wbs_dat_o[29] = net377;
 assign wbs_dat_o[2] = net350;
 assign wbs_dat_o[30] = net378;
 assign wbs_dat_o[31] = net379;
 assign wbs_dat_o[3] = net351;
 assign wbs_dat_o[4] = net352;
 assign wbs_dat_o[5] = net353;
 assign wbs_dat_o[6] = net354;
 assign wbs_dat_o[7] = net355;
 assign wbs_dat_o[8] = net356;
 assign wbs_dat_o[9] = net357;
endmodule

