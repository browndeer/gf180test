VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 680.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 443.520 4.000 444.080 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 450.240 4.000 450.800 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 386.400 4.000 386.960 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 262.080 4.000 262.640 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 225.120 4.000 225.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 676.000 299.600 679.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 168.000 599.000 168.560 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 641.760 599.000 642.320 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 676.000 390.320 679.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 26.880 599.000 27.440 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 676.000 37.520 679.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 676.000 470.960 679.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 1.000 450.800 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 676.000 598.640 679.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 594.720 599.000 595.280 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1.000 528.080 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 534.240 4.000 534.800 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 436.800 4.000 437.360 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 497.280 4.000 497.840 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 675.360 599.000 675.920 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 1.000 417.200 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.800 4.000 269.360 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 1.000 541.520 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 67.200 4.000 67.760 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 571.200 4.000 571.760 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 676.000 531.440 679.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 604.800 599.000 605.360 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 527.520 599.000 528.080 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 668.640 599.000 669.200 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 329.280 599.000 329.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.960 4.000 121.520 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 161.280 599.000 161.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 676.000 484.400 679.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 295.680 4.000 296.240 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 332.640 4.000 333.200 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 490.560 599.000 491.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 453.600 599.000 454.160 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.640 4.000 165.200 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 1.000 585.200 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 676.000 366.800 679.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 1.000 185.360 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 1.000 61.040 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 672.000 4.000 672.560 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 676.000 185.360 679.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 676.000 131.600 679.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 676.000 329.840 679.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 1.000 548.240 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 204.960 599.000 205.520 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 676.000 581.840 679.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 184.800 4.000 185.360 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.720 4.000 91.280 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 584.640 4.000 585.200 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 1.000 534.800 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 651.840 4.000 652.400 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 366.240 599.000 366.800 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 285.600 599.000 286.160 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 0.000 599.000 0.560 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.880 4.000 195.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 676.000 521.360 679.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 144.480 599.000 145.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 524.160 4.000 524.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 618.240 599.000 618.800 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 676.000 316.400 679.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 299.040 599.000 299.600 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 480.480 4.000 481.040 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 676.000 427.280 679.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 504.000 4.000 504.560 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 676.000 266.000 679.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 319.200 4.000 319.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 661.920 599.000 662.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 676.000 64.400 679.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 676.000 155.120 679.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 1.000 413.840 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 676.000 588.560 679.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 638.400 4.000 638.960 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.760 4.000 474.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1.000 259.280 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 574.560 599.000 575.120 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 1.000 74.480 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1.000 598.640 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 676.000 101.360 679.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 1.000 40.880 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 100.800 599.000 101.360 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 423.360 4.000 423.920 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 181.440 599.000 182.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 238.560 4.000 239.120 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 1.000 561.680 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 57.120 599.000 57.680 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1.000 269.360 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 1.000 215.600 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 676.000 410.480 679.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1.000 437.360 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 265.440 599.000 266.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 676.000 544.880 679.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 1.000 225.680 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 676.000 360.080 679.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 231.840 4.000 232.400 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 1.000 423.920 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 1.000 380.240 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1.000 151.760 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 30.240 4.000 30.800 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 676.000 255.920 679.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 1.000 296.240 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 676.000 229.040 679.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 114.240 4.000 114.800 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 1.000 467.600 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 1.000 165.200 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 325.920 4.000 326.480 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 638.400 599.000 638.960 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 322.560 599.000 323.120 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1.000 195.440 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 676.000 218.960 679.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 561.120 4.000 561.680 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 500.640 599.000 501.200 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 676.000 20.720 679.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 137.760 599.000 138.320 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 676.000 279.440 679.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.440 4.000 98.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 676.000 108.080 679.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 174.720 599.000 175.280 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 487.200 4.000 487.760 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 282.240 4.000 282.800 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 520.800 599.000 521.360 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 676.000 286.160 679.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 676.000 94.640 679.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 676.000 353.360 679.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 577.920 4.000 578.480 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 601.440 4.000 602.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 198.240 599.000 198.800 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 676.000 242.480 679.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 47.040 4.000 47.600 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 676.000 501.200 679.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.720 4.000 259.280 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 430.080 4.000 430.640 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 676.000 7.280 679.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 564.480 4.000 565.040 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 1.000 454.160 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 628.320 4.000 628.880 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1.000 289.520 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 676.000 309.680 679.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 389.760 599.000 390.320 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 1.000 306.320 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 215.040 4.000 215.600 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 676.000 561.680 679.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 43.680 599.000 44.240 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 1.000 208.880 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 507.360 599.000 507.920 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 676.000 259.280 679.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 676.000 205.520 679.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 676.000 14.000 679.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 676.000 212.240 679.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 1.000 299.600 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 255.360 599.000 255.920 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 676.000 457.520 679.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 676.000 413.840 679.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.360 4.000 171.920 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 188.160 4.000 188.720 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 658.560 4.000 659.120 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 1.000 232.400 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 624.960 599.000 625.520 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 1.000 111.440 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 463.680 599.000 464.240 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.800 4.000 17.360 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 1.000 376.880 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 676.000 124.880 679.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 1.000 128.240 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 272.160 599.000 272.720 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 10.080 4.000 10.640 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 676.000 538.160 679.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 676.000 514.640 679.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 383.040 599.000 383.600 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 23.520 4.000 24.080 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 460.320 4.000 460.880 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 1.000 239.120 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 302.400 599.000 302.960 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 547.680 4.000 548.240 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 396.480 599.000 397.040 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 676.000 272.720 679.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 567.840 599.000 568.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 1.000 339.920 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 339.360 599.000 339.920 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 131.040 599.000 131.600 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 635.040 4.000 635.600 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 440.160 599.000 440.720 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 1.000 188.720 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.960 4.000 289.520 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 1.000 343.280 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 621.600 4.000 622.160 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 676.000 346.640 679.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 551.040 599.000 551.600 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 1.000 276.080 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 147.840 4.000 148.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 336.000 599.000 336.560 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 70.560 599.000 71.120 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 676.000 336.560 679.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 154.560 599.000 155.120 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 1.000 313.040 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 676.000 302.960 679.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 557.760 599.000 558.320 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 292.320 599.000 292.880 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 50.400 599.000 50.960 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 124.320 599.000 124.880 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 104.160 4.000 104.720 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 20.160 599.000 20.720 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 235.200 599.000 235.760 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 581.280 599.000 581.840 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 1.000 37.520 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1.000 262.640 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 676.000 57.680 679.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 676.000 50.960 679.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 453.600 4.000 454.160 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 1.000 148.400 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 1.000 578.480 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 676.000 323.120 679.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 676.000 182.000 679.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 614.880 4.000 615.440 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 80.640 599.000 81.200 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 608.160 4.000 608.720 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 477.120 599.000 477.680 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 676.000 198.800 679.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 191.520 599.000 192.080 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 676.000 447.440 679.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 483.840 599.000 484.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 245.280 4.000 245.840 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 420.000 599.000 420.560 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 676.000 477.680 679.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1.000 171.920 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 1.000 554.960 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 87.360 599.000 87.920 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 225.120 599.000 225.680 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 676.000 575.120 679.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 36.960 4.000 37.520 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 346.080 599.000 346.640 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 278.880 599.000 279.440 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 493.920 599.000 494.480 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 403.200 599.000 403.760 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 645.120 4.000 645.680 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 510.720 4.000 511.280 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1.000 474.320 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1.000 565.040 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 1.000 91.280 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.280 4.000 77.840 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 676.000 0.560 679.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 94.080 599.000 94.640 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 676.000 81.200 679.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 376.320 4.000 376.880 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 676.000 222.320 679.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 676.000 434.000 679.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 1.000 178.640 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 433.440 599.000 434.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1.000 571.760 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 676.000 87.920 679.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1.000 114.800 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 648.480 599.000 649.040 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 676.000 595.280 679.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 588.000 599.000 588.560 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 676.000 235.760 679.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 564.480 599.000 565.040 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 1.000 326.480 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 676.000 71.120 679.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1.000 17.360 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 1.000 3.920 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 676.000 44.240 679.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 1.000 333.200 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.520 4.000 276.080 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 349.440 4.000 350.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 117.600 599.000 118.160 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 676.000 192.080 679.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 406.560 4.000 407.120 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 1.000 121.520 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1.000 282.800 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 676.000 487.760 679.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1.000 511.280 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.920 4.000 74.480 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 467.040 4.000 467.600 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 3.360 4.000 3.920 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 598.080 4.000 598.640 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1.000 491.120 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 676.000 168.560 679.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 33.600 599.000 34.160 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 446.880 599.000 447.440 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 342.720 4.000 343.280 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 372.960 599.000 373.520 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 1.000 487.760 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 676.000 524.720 679.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 107.520 599.000 108.080 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 676.000 339.920 679.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 1.000 591.920 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 312.480 4.000 313.040 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 1.000 77.840 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 359.520 599.000 360.080 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 151.200 4.000 151.760 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 456.960 599.000 457.520 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 1.000 158.480 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 6.720 599.000 7.280 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 676.000 145.040 679.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 676.000 507.920 679.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 530.880 599.000 531.440 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 676.000 118.160 679.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 413.280 4.000 413.840 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 662.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 662.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 662.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 662.780 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 662.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 662.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 662.780 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 662.780 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 151.200 599.000 151.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 676.000 74.480 679.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 262.080 599.000 262.640 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 676.000 383.600 679.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 676.000 249.200 679.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 369.600 4.000 370.160 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1.000 54.320 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.480 4.000 61.040 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 470.400 599.000 470.960 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 1.000 407.120 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 241.920 599.000 242.480 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 13.440 599.000 14.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.320 4.000 40.880 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 676.000 558.320 679.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1.000 518.000 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 188.160 599.000 188.720 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 676.000 34.160 679.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 110.880 4.000 111.440 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 1.000 67.760 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 676.000 175.280 679.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 416.640 599.000 417.200 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 655.200 599.000 655.760 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 1.000 252.560 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 252.000 4.000 252.560 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 309.120 599.000 309.680 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 1.000 497.840 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 676.000 450.800 679.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 1.000 481.040 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 157.920 4.000 158.480 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 1.000 30.800 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 40.320 599.000 40.880 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 211.680 599.000 212.240 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 676.000 161.840 679.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 601.440 599.000 602.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.560 4.000 491.120 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 540.960 4.000 541.520 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 517.440 4.000 518.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 1.000 24.080 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.400 4.000 134.960 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 379.680 599.000 380.240 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 1.000 370.160 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 676.000 397.040 679.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 676.000 551.600 679.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1.000 98.000 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 299.040 4.000 299.600 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 676.000 568.400 679.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 379.680 4.000 380.240 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 544.320 599.000 544.880 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 248.640 599.000 249.200 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 1.000 444.080 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 676.000 494.480 679.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 676.000 111.440 679.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 1.000 202.160 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 426.720 599.000 427.280 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 1.000 524.720 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 228.480 599.000 229.040 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 339.360 4.000 339.920 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 63.840 599.000 64.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 1.000 104.720 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 1.000 319.760 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 315.840 599.000 316.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 676.000 464.240 679.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 611.520 599.000 612.080 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 77.280 599.000 77.840 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 127.680 4.000 128.240 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 409.920 599.000 410.480 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 1.000 10.640 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 631.680 599.000 632.240 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 676.000 440.720 679.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 114.240 599.000 114.800 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 676.000 420.560 679.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 178.080 4.000 178.640 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.600 4.000 202.160 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 1.000 430.640 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 1.000 504.560 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 305.760 4.000 306.320 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 554.400 4.000 554.960 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 676.000 138.320 679.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.320 4.000 208.880 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1.000 134.960 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 1.000 47.600 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 676.000 292.880 679.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 676.000 148.400 679.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1.000 350.000 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 676.000 403.760 679.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 218.400 599.000 218.960 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 416.640 4.000 417.200 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 537.600 599.000 538.160 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 1.000 141.680 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 1.000 245.840 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.760 4.000 54.320 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 514.080 599.000 514.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1.000 386.960 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 676.000 376.880 679.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 676.000 373.520 679.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 591.360 4.000 591.920 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 676.000 27.440 679.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 1.000 460.880 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 141.120 4.000 141.680 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.520 4.000 528.080 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 352.800 599.000 353.360 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 593.040 663.450 ;
      LAYER Metal2 ;
        RECT 0.140 679.300 598.500 679.700 ;
        RECT 0.860 675.700 6.420 679.300 ;
        RECT 7.580 675.700 13.140 679.300 ;
        RECT 14.300 675.700 19.860 679.300 ;
        RECT 21.020 675.700 26.580 679.300 ;
        RECT 27.740 675.700 33.300 679.300 ;
        RECT 34.460 675.700 36.660 679.300 ;
        RECT 37.820 675.700 43.380 679.300 ;
        RECT 44.540 675.700 50.100 679.300 ;
        RECT 51.260 675.700 56.820 679.300 ;
        RECT 57.980 675.700 63.540 679.300 ;
        RECT 64.700 675.700 70.260 679.300 ;
        RECT 71.420 675.700 73.620 679.300 ;
        RECT 74.780 675.700 80.340 679.300 ;
        RECT 81.500 675.700 87.060 679.300 ;
        RECT 88.220 675.700 93.780 679.300 ;
        RECT 94.940 675.700 100.500 679.300 ;
        RECT 101.660 675.700 107.220 679.300 ;
        RECT 108.380 675.700 110.580 679.300 ;
        RECT 111.740 675.700 117.300 679.300 ;
        RECT 118.460 675.700 124.020 679.300 ;
        RECT 125.180 675.700 130.740 679.300 ;
        RECT 131.900 675.700 137.460 679.300 ;
        RECT 138.620 675.700 144.180 679.300 ;
        RECT 145.340 675.700 147.540 679.300 ;
        RECT 148.700 675.700 154.260 679.300 ;
        RECT 155.420 675.700 160.980 679.300 ;
        RECT 162.140 675.700 167.700 679.300 ;
        RECT 168.860 675.700 174.420 679.300 ;
        RECT 175.580 675.700 181.140 679.300 ;
        RECT 182.300 675.700 184.500 679.300 ;
        RECT 185.660 675.700 191.220 679.300 ;
        RECT 192.380 675.700 197.940 679.300 ;
        RECT 199.100 675.700 204.660 679.300 ;
        RECT 205.820 675.700 211.380 679.300 ;
        RECT 212.540 675.700 218.100 679.300 ;
        RECT 219.260 675.700 221.460 679.300 ;
        RECT 222.620 675.700 228.180 679.300 ;
        RECT 229.340 675.700 234.900 679.300 ;
        RECT 236.060 675.700 241.620 679.300 ;
        RECT 242.780 675.700 248.340 679.300 ;
        RECT 249.500 675.700 255.060 679.300 ;
        RECT 256.220 675.700 258.420 679.300 ;
        RECT 259.580 675.700 265.140 679.300 ;
        RECT 266.300 675.700 271.860 679.300 ;
        RECT 273.020 675.700 278.580 679.300 ;
        RECT 279.740 675.700 285.300 679.300 ;
        RECT 286.460 675.700 292.020 679.300 ;
        RECT 293.180 675.700 298.740 679.300 ;
        RECT 299.900 675.700 302.100 679.300 ;
        RECT 303.260 675.700 308.820 679.300 ;
        RECT 309.980 675.700 315.540 679.300 ;
        RECT 316.700 675.700 322.260 679.300 ;
        RECT 323.420 675.700 328.980 679.300 ;
        RECT 330.140 675.700 335.700 679.300 ;
        RECT 336.860 675.700 339.060 679.300 ;
        RECT 340.220 675.700 345.780 679.300 ;
        RECT 346.940 675.700 352.500 679.300 ;
        RECT 353.660 675.700 359.220 679.300 ;
        RECT 360.380 675.700 365.940 679.300 ;
        RECT 367.100 675.700 372.660 679.300 ;
        RECT 373.820 675.700 376.020 679.300 ;
        RECT 377.180 675.700 382.740 679.300 ;
        RECT 383.900 675.700 389.460 679.300 ;
        RECT 390.620 675.700 396.180 679.300 ;
        RECT 397.340 675.700 402.900 679.300 ;
        RECT 404.060 675.700 409.620 679.300 ;
        RECT 410.780 675.700 412.980 679.300 ;
        RECT 414.140 675.700 419.700 679.300 ;
        RECT 420.860 675.700 426.420 679.300 ;
        RECT 427.580 675.700 433.140 679.300 ;
        RECT 434.300 675.700 439.860 679.300 ;
        RECT 441.020 675.700 446.580 679.300 ;
        RECT 447.740 675.700 449.940 679.300 ;
        RECT 451.100 675.700 456.660 679.300 ;
        RECT 457.820 675.700 463.380 679.300 ;
        RECT 464.540 675.700 470.100 679.300 ;
        RECT 471.260 675.700 476.820 679.300 ;
        RECT 477.980 675.700 483.540 679.300 ;
        RECT 484.700 675.700 486.900 679.300 ;
        RECT 488.060 675.700 493.620 679.300 ;
        RECT 494.780 675.700 500.340 679.300 ;
        RECT 501.500 675.700 507.060 679.300 ;
        RECT 508.220 675.700 513.780 679.300 ;
        RECT 514.940 675.700 520.500 679.300 ;
        RECT 521.660 675.700 523.860 679.300 ;
        RECT 525.020 675.700 530.580 679.300 ;
        RECT 531.740 675.700 537.300 679.300 ;
        RECT 538.460 675.700 544.020 679.300 ;
        RECT 545.180 675.700 550.740 679.300 ;
        RECT 551.900 675.700 557.460 679.300 ;
        RECT 558.620 675.700 560.820 679.300 ;
        RECT 561.980 675.700 567.540 679.300 ;
        RECT 568.700 675.700 574.260 679.300 ;
        RECT 575.420 675.700 580.980 679.300 ;
        RECT 582.140 675.700 587.700 679.300 ;
        RECT 588.860 675.700 594.420 679.300 ;
        RECT 595.580 675.700 597.780 679.300 ;
        RECT 0.140 4.300 598.500 675.700 ;
        RECT 0.860 0.700 3.060 4.300 ;
        RECT 4.220 0.700 9.780 4.300 ;
        RECT 10.940 0.700 16.500 4.300 ;
        RECT 17.660 0.700 23.220 4.300 ;
        RECT 24.380 0.700 29.940 4.300 ;
        RECT 31.100 0.700 36.660 4.300 ;
        RECT 37.820 0.700 40.020 4.300 ;
        RECT 41.180 0.700 46.740 4.300 ;
        RECT 47.900 0.700 53.460 4.300 ;
        RECT 54.620 0.700 60.180 4.300 ;
        RECT 61.340 0.700 66.900 4.300 ;
        RECT 68.060 0.700 73.620 4.300 ;
        RECT 74.780 0.700 76.980 4.300 ;
        RECT 78.140 0.700 83.700 4.300 ;
        RECT 84.860 0.700 90.420 4.300 ;
        RECT 91.580 0.700 97.140 4.300 ;
        RECT 98.300 0.700 103.860 4.300 ;
        RECT 105.020 0.700 110.580 4.300 ;
        RECT 111.740 0.700 113.940 4.300 ;
        RECT 115.100 0.700 120.660 4.300 ;
        RECT 121.820 0.700 127.380 4.300 ;
        RECT 128.540 0.700 134.100 4.300 ;
        RECT 135.260 0.700 140.820 4.300 ;
        RECT 141.980 0.700 147.540 4.300 ;
        RECT 148.700 0.700 150.900 4.300 ;
        RECT 152.060 0.700 157.620 4.300 ;
        RECT 158.780 0.700 164.340 4.300 ;
        RECT 165.500 0.700 171.060 4.300 ;
        RECT 172.220 0.700 177.780 4.300 ;
        RECT 178.940 0.700 184.500 4.300 ;
        RECT 185.660 0.700 187.860 4.300 ;
        RECT 189.020 0.700 194.580 4.300 ;
        RECT 195.740 0.700 201.300 4.300 ;
        RECT 202.460 0.700 208.020 4.300 ;
        RECT 209.180 0.700 214.740 4.300 ;
        RECT 215.900 0.700 221.460 4.300 ;
        RECT 222.620 0.700 224.820 4.300 ;
        RECT 225.980 0.700 231.540 4.300 ;
        RECT 232.700 0.700 238.260 4.300 ;
        RECT 239.420 0.700 244.980 4.300 ;
        RECT 246.140 0.700 251.700 4.300 ;
        RECT 252.860 0.700 258.420 4.300 ;
        RECT 259.580 0.700 261.780 4.300 ;
        RECT 262.940 0.700 268.500 4.300 ;
        RECT 269.660 0.700 275.220 4.300 ;
        RECT 276.380 0.700 281.940 4.300 ;
        RECT 283.100 0.700 288.660 4.300 ;
        RECT 289.820 0.700 295.380 4.300 ;
        RECT 296.540 0.700 298.740 4.300 ;
        RECT 299.900 0.700 305.460 4.300 ;
        RECT 306.620 0.700 312.180 4.300 ;
        RECT 313.340 0.700 318.900 4.300 ;
        RECT 320.060 0.700 325.620 4.300 ;
        RECT 326.780 0.700 332.340 4.300 ;
        RECT 333.500 0.700 339.060 4.300 ;
        RECT 340.220 0.700 342.420 4.300 ;
        RECT 343.580 0.700 349.140 4.300 ;
        RECT 350.300 0.700 355.860 4.300 ;
        RECT 357.020 0.700 362.580 4.300 ;
        RECT 363.740 0.700 369.300 4.300 ;
        RECT 370.460 0.700 376.020 4.300 ;
        RECT 377.180 0.700 379.380 4.300 ;
        RECT 380.540 0.700 386.100 4.300 ;
        RECT 387.260 0.700 392.820 4.300 ;
        RECT 393.980 0.700 399.540 4.300 ;
        RECT 400.700 0.700 406.260 4.300 ;
        RECT 407.420 0.700 412.980 4.300 ;
        RECT 414.140 0.700 416.340 4.300 ;
        RECT 417.500 0.700 423.060 4.300 ;
        RECT 424.220 0.700 429.780 4.300 ;
        RECT 430.940 0.700 436.500 4.300 ;
        RECT 437.660 0.700 443.220 4.300 ;
        RECT 444.380 0.700 449.940 4.300 ;
        RECT 451.100 0.700 453.300 4.300 ;
        RECT 454.460 0.700 460.020 4.300 ;
        RECT 461.180 0.700 466.740 4.300 ;
        RECT 467.900 0.700 473.460 4.300 ;
        RECT 474.620 0.700 480.180 4.300 ;
        RECT 481.340 0.700 486.900 4.300 ;
        RECT 488.060 0.700 490.260 4.300 ;
        RECT 491.420 0.700 496.980 4.300 ;
        RECT 498.140 0.700 503.700 4.300 ;
        RECT 504.860 0.700 510.420 4.300 ;
        RECT 511.580 0.700 517.140 4.300 ;
        RECT 518.300 0.700 523.860 4.300 ;
        RECT 525.020 0.700 527.220 4.300 ;
        RECT 528.380 0.700 533.940 4.300 ;
        RECT 535.100 0.700 540.660 4.300 ;
        RECT 541.820 0.700 547.380 4.300 ;
        RECT 548.540 0.700 554.100 4.300 ;
        RECT 555.260 0.700 560.820 4.300 ;
        RECT 561.980 0.700 564.180 4.300 ;
        RECT 565.340 0.700 570.900 4.300 ;
        RECT 572.060 0.700 577.620 4.300 ;
        RECT 578.780 0.700 584.340 4.300 ;
        RECT 585.500 0.700 591.060 4.300 ;
        RECT 592.220 0.700 597.780 4.300 ;
        RECT 0.140 0.090 598.500 0.700 ;
      LAYER Metal3 ;
        RECT 0.090 675.060 595.700 675.780 ;
        RECT 0.090 672.860 598.550 675.060 ;
        RECT 0.090 671.700 0.700 672.860 ;
        RECT 4.300 671.700 598.550 672.860 ;
        RECT 0.090 669.500 598.550 671.700 ;
        RECT 0.090 668.340 595.700 669.500 ;
        RECT 0.090 666.140 598.550 668.340 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 598.550 666.140 ;
        RECT 0.090 662.780 598.550 664.980 ;
        RECT 0.090 661.620 595.700 662.780 ;
        RECT 0.090 659.420 598.550 661.620 ;
        RECT 0.090 658.260 0.700 659.420 ;
        RECT 4.300 658.260 598.550 659.420 ;
        RECT 0.090 656.060 598.550 658.260 ;
        RECT 0.090 654.900 595.700 656.060 ;
        RECT 0.090 652.700 598.550 654.900 ;
        RECT 0.090 651.540 0.700 652.700 ;
        RECT 4.300 651.540 598.550 652.700 ;
        RECT 0.090 649.340 598.550 651.540 ;
        RECT 0.090 648.180 595.700 649.340 ;
        RECT 0.090 645.980 598.550 648.180 ;
        RECT 0.090 644.820 0.700 645.980 ;
        RECT 4.300 644.820 598.550 645.980 ;
        RECT 0.090 642.620 598.550 644.820 ;
        RECT 0.090 641.460 595.700 642.620 ;
        RECT 0.090 639.260 598.550 641.460 ;
        RECT 0.090 638.100 0.700 639.260 ;
        RECT 4.300 638.100 595.700 639.260 ;
        RECT 0.090 635.900 598.550 638.100 ;
        RECT 0.090 634.740 0.700 635.900 ;
        RECT 4.300 634.740 598.550 635.900 ;
        RECT 0.090 632.540 598.550 634.740 ;
        RECT 0.090 631.380 595.700 632.540 ;
        RECT 0.090 629.180 598.550 631.380 ;
        RECT 0.090 628.020 0.700 629.180 ;
        RECT 4.300 628.020 598.550 629.180 ;
        RECT 0.090 625.820 598.550 628.020 ;
        RECT 0.090 624.660 595.700 625.820 ;
        RECT 0.090 622.460 598.550 624.660 ;
        RECT 0.090 621.300 0.700 622.460 ;
        RECT 4.300 621.300 598.550 622.460 ;
        RECT 0.090 619.100 598.550 621.300 ;
        RECT 0.090 617.940 595.700 619.100 ;
        RECT 0.090 615.740 598.550 617.940 ;
        RECT 0.090 614.580 0.700 615.740 ;
        RECT 4.300 614.580 598.550 615.740 ;
        RECT 0.090 612.380 598.550 614.580 ;
        RECT 0.090 611.220 595.700 612.380 ;
        RECT 0.090 609.020 598.550 611.220 ;
        RECT 0.090 607.860 0.700 609.020 ;
        RECT 4.300 607.860 598.550 609.020 ;
        RECT 0.090 605.660 598.550 607.860 ;
        RECT 0.090 604.500 595.700 605.660 ;
        RECT 0.090 602.300 598.550 604.500 ;
        RECT 0.090 601.140 0.700 602.300 ;
        RECT 4.300 601.140 595.700 602.300 ;
        RECT 0.090 598.940 598.550 601.140 ;
        RECT 0.090 597.780 0.700 598.940 ;
        RECT 4.300 597.780 598.550 598.940 ;
        RECT 0.090 595.580 598.550 597.780 ;
        RECT 0.090 594.420 595.700 595.580 ;
        RECT 0.090 592.220 598.550 594.420 ;
        RECT 0.090 591.060 0.700 592.220 ;
        RECT 4.300 591.060 598.550 592.220 ;
        RECT 0.090 588.860 598.550 591.060 ;
        RECT 0.090 587.700 595.700 588.860 ;
        RECT 0.090 585.500 598.550 587.700 ;
        RECT 0.090 584.340 0.700 585.500 ;
        RECT 4.300 584.340 598.550 585.500 ;
        RECT 0.090 582.140 598.550 584.340 ;
        RECT 0.090 580.980 595.700 582.140 ;
        RECT 0.090 578.780 598.550 580.980 ;
        RECT 0.090 577.620 0.700 578.780 ;
        RECT 4.300 577.620 598.550 578.780 ;
        RECT 0.090 575.420 598.550 577.620 ;
        RECT 0.090 574.260 595.700 575.420 ;
        RECT 0.090 572.060 598.550 574.260 ;
        RECT 0.090 570.900 0.700 572.060 ;
        RECT 4.300 570.900 598.550 572.060 ;
        RECT 0.090 568.700 598.550 570.900 ;
        RECT 0.090 567.540 595.700 568.700 ;
        RECT 0.090 565.340 598.550 567.540 ;
        RECT 0.090 564.180 0.700 565.340 ;
        RECT 4.300 564.180 595.700 565.340 ;
        RECT 0.090 561.980 598.550 564.180 ;
        RECT 0.090 560.820 0.700 561.980 ;
        RECT 4.300 560.820 598.550 561.980 ;
        RECT 0.090 558.620 598.550 560.820 ;
        RECT 0.090 557.460 595.700 558.620 ;
        RECT 0.090 555.260 598.550 557.460 ;
        RECT 0.090 554.100 0.700 555.260 ;
        RECT 4.300 554.100 598.550 555.260 ;
        RECT 0.090 551.900 598.550 554.100 ;
        RECT 0.090 550.740 595.700 551.900 ;
        RECT 0.090 548.540 598.550 550.740 ;
        RECT 0.090 547.380 0.700 548.540 ;
        RECT 4.300 547.380 598.550 548.540 ;
        RECT 0.090 545.180 598.550 547.380 ;
        RECT 0.090 544.020 595.700 545.180 ;
        RECT 0.090 541.820 598.550 544.020 ;
        RECT 0.090 540.660 0.700 541.820 ;
        RECT 4.300 540.660 598.550 541.820 ;
        RECT 0.090 538.460 598.550 540.660 ;
        RECT 0.090 537.300 595.700 538.460 ;
        RECT 0.090 535.100 598.550 537.300 ;
        RECT 0.090 533.940 0.700 535.100 ;
        RECT 4.300 533.940 598.550 535.100 ;
        RECT 0.090 531.740 598.550 533.940 ;
        RECT 0.090 530.580 595.700 531.740 ;
        RECT 0.090 528.380 598.550 530.580 ;
        RECT 0.090 527.220 0.700 528.380 ;
        RECT 4.300 527.220 595.700 528.380 ;
        RECT 0.090 525.020 598.550 527.220 ;
        RECT 0.090 523.860 0.700 525.020 ;
        RECT 4.300 523.860 598.550 525.020 ;
        RECT 0.090 521.660 598.550 523.860 ;
        RECT 0.090 520.500 595.700 521.660 ;
        RECT 0.090 518.300 598.550 520.500 ;
        RECT 0.090 517.140 0.700 518.300 ;
        RECT 4.300 517.140 598.550 518.300 ;
        RECT 0.090 514.940 598.550 517.140 ;
        RECT 0.090 513.780 595.700 514.940 ;
        RECT 0.090 511.580 598.550 513.780 ;
        RECT 0.090 510.420 0.700 511.580 ;
        RECT 4.300 510.420 598.550 511.580 ;
        RECT 0.090 508.220 598.550 510.420 ;
        RECT 0.090 507.060 595.700 508.220 ;
        RECT 0.090 504.860 598.550 507.060 ;
        RECT 0.090 503.700 0.700 504.860 ;
        RECT 4.300 503.700 598.550 504.860 ;
        RECT 0.090 501.500 598.550 503.700 ;
        RECT 0.090 500.340 595.700 501.500 ;
        RECT 0.090 498.140 598.550 500.340 ;
        RECT 0.090 496.980 0.700 498.140 ;
        RECT 4.300 496.980 598.550 498.140 ;
        RECT 0.090 494.780 598.550 496.980 ;
        RECT 0.090 493.620 595.700 494.780 ;
        RECT 0.090 491.420 598.550 493.620 ;
        RECT 0.090 490.260 0.700 491.420 ;
        RECT 4.300 490.260 595.700 491.420 ;
        RECT 0.090 488.060 598.550 490.260 ;
        RECT 0.090 486.900 0.700 488.060 ;
        RECT 4.300 486.900 598.550 488.060 ;
        RECT 0.090 484.700 598.550 486.900 ;
        RECT 0.090 483.540 595.700 484.700 ;
        RECT 0.090 481.340 598.550 483.540 ;
        RECT 0.090 480.180 0.700 481.340 ;
        RECT 4.300 480.180 598.550 481.340 ;
        RECT 0.090 477.980 598.550 480.180 ;
        RECT 0.090 476.820 595.700 477.980 ;
        RECT 0.090 474.620 598.550 476.820 ;
        RECT 0.090 473.460 0.700 474.620 ;
        RECT 4.300 473.460 598.550 474.620 ;
        RECT 0.090 471.260 598.550 473.460 ;
        RECT 0.090 470.100 595.700 471.260 ;
        RECT 0.090 467.900 598.550 470.100 ;
        RECT 0.090 466.740 0.700 467.900 ;
        RECT 4.300 466.740 598.550 467.900 ;
        RECT 0.090 464.540 598.550 466.740 ;
        RECT 0.090 463.380 595.700 464.540 ;
        RECT 0.090 461.180 598.550 463.380 ;
        RECT 0.090 460.020 0.700 461.180 ;
        RECT 4.300 460.020 598.550 461.180 ;
        RECT 0.090 457.820 598.550 460.020 ;
        RECT 0.090 456.660 595.700 457.820 ;
        RECT 0.090 454.460 598.550 456.660 ;
        RECT 0.090 453.300 0.700 454.460 ;
        RECT 4.300 453.300 595.700 454.460 ;
        RECT 0.090 451.100 598.550 453.300 ;
        RECT 0.090 449.940 0.700 451.100 ;
        RECT 4.300 449.940 598.550 451.100 ;
        RECT 0.090 447.740 598.550 449.940 ;
        RECT 0.090 446.580 595.700 447.740 ;
        RECT 0.090 444.380 598.550 446.580 ;
        RECT 0.090 443.220 0.700 444.380 ;
        RECT 4.300 443.220 598.550 444.380 ;
        RECT 0.090 441.020 598.550 443.220 ;
        RECT 0.090 439.860 595.700 441.020 ;
        RECT 0.090 437.660 598.550 439.860 ;
        RECT 0.090 436.500 0.700 437.660 ;
        RECT 4.300 436.500 598.550 437.660 ;
        RECT 0.090 434.300 598.550 436.500 ;
        RECT 0.090 433.140 595.700 434.300 ;
        RECT 0.090 430.940 598.550 433.140 ;
        RECT 0.090 429.780 0.700 430.940 ;
        RECT 4.300 429.780 598.550 430.940 ;
        RECT 0.090 427.580 598.550 429.780 ;
        RECT 0.090 426.420 595.700 427.580 ;
        RECT 0.090 424.220 598.550 426.420 ;
        RECT 0.090 423.060 0.700 424.220 ;
        RECT 4.300 423.060 598.550 424.220 ;
        RECT 0.090 420.860 598.550 423.060 ;
        RECT 0.090 419.700 595.700 420.860 ;
        RECT 0.090 417.500 598.550 419.700 ;
        RECT 0.090 416.340 0.700 417.500 ;
        RECT 4.300 416.340 595.700 417.500 ;
        RECT 0.090 414.140 598.550 416.340 ;
        RECT 0.090 412.980 0.700 414.140 ;
        RECT 4.300 412.980 598.550 414.140 ;
        RECT 0.090 410.780 598.550 412.980 ;
        RECT 0.090 409.620 595.700 410.780 ;
        RECT 0.090 407.420 598.550 409.620 ;
        RECT 0.090 406.260 0.700 407.420 ;
        RECT 4.300 406.260 598.550 407.420 ;
        RECT 0.090 404.060 598.550 406.260 ;
        RECT 0.090 402.900 595.700 404.060 ;
        RECT 0.090 400.700 598.550 402.900 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 598.550 400.700 ;
        RECT 0.090 397.340 598.550 399.540 ;
        RECT 0.090 396.180 595.700 397.340 ;
        RECT 0.090 393.980 598.550 396.180 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 598.550 393.980 ;
        RECT 0.090 390.620 598.550 392.820 ;
        RECT 0.090 389.460 595.700 390.620 ;
        RECT 0.090 387.260 598.550 389.460 ;
        RECT 0.090 386.100 0.700 387.260 ;
        RECT 4.300 386.100 598.550 387.260 ;
        RECT 0.090 383.900 598.550 386.100 ;
        RECT 0.090 382.740 595.700 383.900 ;
        RECT 0.090 380.540 598.550 382.740 ;
        RECT 0.090 379.380 0.700 380.540 ;
        RECT 4.300 379.380 595.700 380.540 ;
        RECT 0.090 377.180 598.550 379.380 ;
        RECT 0.090 376.020 0.700 377.180 ;
        RECT 4.300 376.020 598.550 377.180 ;
        RECT 0.090 373.820 598.550 376.020 ;
        RECT 0.090 372.660 595.700 373.820 ;
        RECT 0.090 370.460 598.550 372.660 ;
        RECT 0.090 369.300 0.700 370.460 ;
        RECT 4.300 369.300 598.550 370.460 ;
        RECT 0.090 367.100 598.550 369.300 ;
        RECT 0.090 365.940 595.700 367.100 ;
        RECT 0.090 363.740 598.550 365.940 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 598.550 363.740 ;
        RECT 0.090 360.380 598.550 362.580 ;
        RECT 0.090 359.220 595.700 360.380 ;
        RECT 0.090 357.020 598.550 359.220 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 598.550 357.020 ;
        RECT 0.090 353.660 598.550 355.860 ;
        RECT 0.090 352.500 595.700 353.660 ;
        RECT 0.090 350.300 598.550 352.500 ;
        RECT 0.090 349.140 0.700 350.300 ;
        RECT 4.300 349.140 598.550 350.300 ;
        RECT 0.090 346.940 598.550 349.140 ;
        RECT 0.090 345.780 595.700 346.940 ;
        RECT 0.090 343.580 598.550 345.780 ;
        RECT 0.090 342.420 0.700 343.580 ;
        RECT 4.300 342.420 598.550 343.580 ;
        RECT 0.090 340.220 598.550 342.420 ;
        RECT 0.090 339.060 0.700 340.220 ;
        RECT 4.300 339.060 595.700 340.220 ;
        RECT 0.090 336.860 598.550 339.060 ;
        RECT 0.090 335.700 595.700 336.860 ;
        RECT 0.090 333.500 598.550 335.700 ;
        RECT 0.090 332.340 0.700 333.500 ;
        RECT 4.300 332.340 598.550 333.500 ;
        RECT 0.090 330.140 598.550 332.340 ;
        RECT 0.090 328.980 595.700 330.140 ;
        RECT 0.090 326.780 598.550 328.980 ;
        RECT 0.090 325.620 0.700 326.780 ;
        RECT 4.300 325.620 598.550 326.780 ;
        RECT 0.090 323.420 598.550 325.620 ;
        RECT 0.090 322.260 595.700 323.420 ;
        RECT 0.090 320.060 598.550 322.260 ;
        RECT 0.090 318.900 0.700 320.060 ;
        RECT 4.300 318.900 598.550 320.060 ;
        RECT 0.090 316.700 598.550 318.900 ;
        RECT 0.090 315.540 595.700 316.700 ;
        RECT 0.090 313.340 598.550 315.540 ;
        RECT 0.090 312.180 0.700 313.340 ;
        RECT 4.300 312.180 598.550 313.340 ;
        RECT 0.090 309.980 598.550 312.180 ;
        RECT 0.090 308.820 595.700 309.980 ;
        RECT 0.090 306.620 598.550 308.820 ;
        RECT 0.090 305.460 0.700 306.620 ;
        RECT 4.300 305.460 598.550 306.620 ;
        RECT 0.090 303.260 598.550 305.460 ;
        RECT 0.090 302.100 595.700 303.260 ;
        RECT 0.090 299.900 598.550 302.100 ;
        RECT 0.090 298.740 0.700 299.900 ;
        RECT 4.300 298.740 595.700 299.900 ;
        RECT 0.090 296.540 598.550 298.740 ;
        RECT 0.090 295.380 0.700 296.540 ;
        RECT 4.300 295.380 598.550 296.540 ;
        RECT 0.090 293.180 598.550 295.380 ;
        RECT 0.090 292.020 595.700 293.180 ;
        RECT 0.090 289.820 598.550 292.020 ;
        RECT 0.090 288.660 0.700 289.820 ;
        RECT 4.300 288.660 598.550 289.820 ;
        RECT 0.090 286.460 598.550 288.660 ;
        RECT 0.090 285.300 595.700 286.460 ;
        RECT 0.090 283.100 598.550 285.300 ;
        RECT 0.090 281.940 0.700 283.100 ;
        RECT 4.300 281.940 598.550 283.100 ;
        RECT 0.090 279.740 598.550 281.940 ;
        RECT 0.090 278.580 595.700 279.740 ;
        RECT 0.090 276.380 598.550 278.580 ;
        RECT 0.090 275.220 0.700 276.380 ;
        RECT 4.300 275.220 598.550 276.380 ;
        RECT 0.090 273.020 598.550 275.220 ;
        RECT 0.090 271.860 595.700 273.020 ;
        RECT 0.090 269.660 598.550 271.860 ;
        RECT 0.090 268.500 0.700 269.660 ;
        RECT 4.300 268.500 598.550 269.660 ;
        RECT 0.090 266.300 598.550 268.500 ;
        RECT 0.090 265.140 595.700 266.300 ;
        RECT 0.090 262.940 598.550 265.140 ;
        RECT 0.090 261.780 0.700 262.940 ;
        RECT 4.300 261.780 595.700 262.940 ;
        RECT 0.090 259.580 598.550 261.780 ;
        RECT 0.090 258.420 0.700 259.580 ;
        RECT 4.300 258.420 598.550 259.580 ;
        RECT 0.090 256.220 598.550 258.420 ;
        RECT 0.090 255.060 595.700 256.220 ;
        RECT 0.090 252.860 598.550 255.060 ;
        RECT 0.090 251.700 0.700 252.860 ;
        RECT 4.300 251.700 598.550 252.860 ;
        RECT 0.090 249.500 598.550 251.700 ;
        RECT 0.090 248.340 595.700 249.500 ;
        RECT 0.090 246.140 598.550 248.340 ;
        RECT 0.090 244.980 0.700 246.140 ;
        RECT 4.300 244.980 598.550 246.140 ;
        RECT 0.090 242.780 598.550 244.980 ;
        RECT 0.090 241.620 595.700 242.780 ;
        RECT 0.090 239.420 598.550 241.620 ;
        RECT 0.090 238.260 0.700 239.420 ;
        RECT 4.300 238.260 598.550 239.420 ;
        RECT 0.090 236.060 598.550 238.260 ;
        RECT 0.090 234.900 595.700 236.060 ;
        RECT 0.090 232.700 598.550 234.900 ;
        RECT 0.090 231.540 0.700 232.700 ;
        RECT 4.300 231.540 598.550 232.700 ;
        RECT 0.090 229.340 598.550 231.540 ;
        RECT 0.090 228.180 595.700 229.340 ;
        RECT 0.090 225.980 598.550 228.180 ;
        RECT 0.090 224.820 0.700 225.980 ;
        RECT 4.300 224.820 595.700 225.980 ;
        RECT 0.090 222.620 598.550 224.820 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 598.550 222.620 ;
        RECT 0.090 219.260 598.550 221.460 ;
        RECT 0.090 218.100 595.700 219.260 ;
        RECT 0.090 215.900 598.550 218.100 ;
        RECT 0.090 214.740 0.700 215.900 ;
        RECT 4.300 214.740 598.550 215.900 ;
        RECT 0.090 212.540 598.550 214.740 ;
        RECT 0.090 211.380 595.700 212.540 ;
        RECT 0.090 209.180 598.550 211.380 ;
        RECT 0.090 208.020 0.700 209.180 ;
        RECT 4.300 208.020 598.550 209.180 ;
        RECT 0.090 205.820 598.550 208.020 ;
        RECT 0.090 204.660 595.700 205.820 ;
        RECT 0.090 202.460 598.550 204.660 ;
        RECT 0.090 201.300 0.700 202.460 ;
        RECT 4.300 201.300 598.550 202.460 ;
        RECT 0.090 199.100 598.550 201.300 ;
        RECT 0.090 197.940 595.700 199.100 ;
        RECT 0.090 195.740 598.550 197.940 ;
        RECT 0.090 194.580 0.700 195.740 ;
        RECT 4.300 194.580 598.550 195.740 ;
        RECT 0.090 192.380 598.550 194.580 ;
        RECT 0.090 191.220 595.700 192.380 ;
        RECT 0.090 189.020 598.550 191.220 ;
        RECT 0.090 187.860 0.700 189.020 ;
        RECT 4.300 187.860 595.700 189.020 ;
        RECT 0.090 185.660 598.550 187.860 ;
        RECT 0.090 184.500 0.700 185.660 ;
        RECT 4.300 184.500 598.550 185.660 ;
        RECT 0.090 182.300 598.550 184.500 ;
        RECT 0.090 181.140 595.700 182.300 ;
        RECT 0.090 178.940 598.550 181.140 ;
        RECT 0.090 177.780 0.700 178.940 ;
        RECT 4.300 177.780 598.550 178.940 ;
        RECT 0.090 175.580 598.550 177.780 ;
        RECT 0.090 174.420 595.700 175.580 ;
        RECT 0.090 172.220 598.550 174.420 ;
        RECT 0.090 171.060 0.700 172.220 ;
        RECT 4.300 171.060 598.550 172.220 ;
        RECT 0.090 168.860 598.550 171.060 ;
        RECT 0.090 167.700 595.700 168.860 ;
        RECT 0.090 165.500 598.550 167.700 ;
        RECT 0.090 164.340 0.700 165.500 ;
        RECT 4.300 164.340 598.550 165.500 ;
        RECT 0.090 162.140 598.550 164.340 ;
        RECT 0.090 160.980 595.700 162.140 ;
        RECT 0.090 158.780 598.550 160.980 ;
        RECT 0.090 157.620 0.700 158.780 ;
        RECT 4.300 157.620 598.550 158.780 ;
        RECT 0.090 155.420 598.550 157.620 ;
        RECT 0.090 154.260 595.700 155.420 ;
        RECT 0.090 152.060 598.550 154.260 ;
        RECT 0.090 150.900 0.700 152.060 ;
        RECT 4.300 150.900 595.700 152.060 ;
        RECT 0.090 148.700 598.550 150.900 ;
        RECT 0.090 147.540 0.700 148.700 ;
        RECT 4.300 147.540 598.550 148.700 ;
        RECT 0.090 145.340 598.550 147.540 ;
        RECT 0.090 144.180 595.700 145.340 ;
        RECT 0.090 141.980 598.550 144.180 ;
        RECT 0.090 140.820 0.700 141.980 ;
        RECT 4.300 140.820 598.550 141.980 ;
        RECT 0.090 138.620 598.550 140.820 ;
        RECT 0.090 137.460 595.700 138.620 ;
        RECT 0.090 135.260 598.550 137.460 ;
        RECT 0.090 134.100 0.700 135.260 ;
        RECT 4.300 134.100 598.550 135.260 ;
        RECT 0.090 131.900 598.550 134.100 ;
        RECT 0.090 130.740 595.700 131.900 ;
        RECT 0.090 128.540 598.550 130.740 ;
        RECT 0.090 127.380 0.700 128.540 ;
        RECT 4.300 127.380 598.550 128.540 ;
        RECT 0.090 125.180 598.550 127.380 ;
        RECT 0.090 124.020 595.700 125.180 ;
        RECT 0.090 121.820 598.550 124.020 ;
        RECT 0.090 120.660 0.700 121.820 ;
        RECT 4.300 120.660 598.550 121.820 ;
        RECT 0.090 118.460 598.550 120.660 ;
        RECT 0.090 117.300 595.700 118.460 ;
        RECT 0.090 115.100 598.550 117.300 ;
        RECT 0.090 113.940 0.700 115.100 ;
        RECT 4.300 113.940 595.700 115.100 ;
        RECT 0.090 111.740 598.550 113.940 ;
        RECT 0.090 110.580 0.700 111.740 ;
        RECT 4.300 110.580 598.550 111.740 ;
        RECT 0.090 108.380 598.550 110.580 ;
        RECT 0.090 107.220 595.700 108.380 ;
        RECT 0.090 105.020 598.550 107.220 ;
        RECT 0.090 103.860 0.700 105.020 ;
        RECT 4.300 103.860 598.550 105.020 ;
        RECT 0.090 101.660 598.550 103.860 ;
        RECT 0.090 100.500 595.700 101.660 ;
        RECT 0.090 98.300 598.550 100.500 ;
        RECT 0.090 97.140 0.700 98.300 ;
        RECT 4.300 97.140 598.550 98.300 ;
        RECT 0.090 94.940 598.550 97.140 ;
        RECT 0.090 93.780 595.700 94.940 ;
        RECT 0.090 91.580 598.550 93.780 ;
        RECT 0.090 90.420 0.700 91.580 ;
        RECT 4.300 90.420 598.550 91.580 ;
        RECT 0.090 88.220 598.550 90.420 ;
        RECT 0.090 87.060 595.700 88.220 ;
        RECT 0.090 84.860 598.550 87.060 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 598.550 84.860 ;
        RECT 0.090 81.500 598.550 83.700 ;
        RECT 0.090 80.340 595.700 81.500 ;
        RECT 0.090 78.140 598.550 80.340 ;
        RECT 0.090 76.980 0.700 78.140 ;
        RECT 4.300 76.980 595.700 78.140 ;
        RECT 0.090 74.780 598.550 76.980 ;
        RECT 0.090 73.620 0.700 74.780 ;
        RECT 4.300 73.620 598.550 74.780 ;
        RECT 0.090 71.420 598.550 73.620 ;
        RECT 0.090 70.260 595.700 71.420 ;
        RECT 0.090 68.060 598.550 70.260 ;
        RECT 0.090 66.900 0.700 68.060 ;
        RECT 4.300 66.900 598.550 68.060 ;
        RECT 0.090 64.700 598.550 66.900 ;
        RECT 0.090 63.540 595.700 64.700 ;
        RECT 0.090 61.340 598.550 63.540 ;
        RECT 0.090 60.180 0.700 61.340 ;
        RECT 4.300 60.180 598.550 61.340 ;
        RECT 0.090 57.980 598.550 60.180 ;
        RECT 0.090 56.820 595.700 57.980 ;
        RECT 0.090 54.620 598.550 56.820 ;
        RECT 0.090 53.460 0.700 54.620 ;
        RECT 4.300 53.460 598.550 54.620 ;
        RECT 0.090 51.260 598.550 53.460 ;
        RECT 0.090 50.100 595.700 51.260 ;
        RECT 0.090 47.900 598.550 50.100 ;
        RECT 0.090 46.740 0.700 47.900 ;
        RECT 4.300 46.740 598.550 47.900 ;
        RECT 0.090 44.540 598.550 46.740 ;
        RECT 0.090 43.380 595.700 44.540 ;
        RECT 0.090 41.180 598.550 43.380 ;
        RECT 0.090 40.020 0.700 41.180 ;
        RECT 4.300 40.020 595.700 41.180 ;
        RECT 0.090 37.820 598.550 40.020 ;
        RECT 0.090 36.660 0.700 37.820 ;
        RECT 4.300 36.660 598.550 37.820 ;
        RECT 0.090 34.460 598.550 36.660 ;
        RECT 0.090 33.300 595.700 34.460 ;
        RECT 0.090 31.100 598.550 33.300 ;
        RECT 0.090 29.940 0.700 31.100 ;
        RECT 4.300 29.940 598.550 31.100 ;
        RECT 0.090 27.740 598.550 29.940 ;
        RECT 0.090 26.580 595.700 27.740 ;
        RECT 0.090 24.380 598.550 26.580 ;
        RECT 0.090 23.220 0.700 24.380 ;
        RECT 4.300 23.220 598.550 24.380 ;
        RECT 0.090 21.020 598.550 23.220 ;
        RECT 0.090 19.860 595.700 21.020 ;
        RECT 0.090 17.660 598.550 19.860 ;
        RECT 0.090 16.500 0.700 17.660 ;
        RECT 4.300 16.500 598.550 17.660 ;
        RECT 0.090 14.300 598.550 16.500 ;
        RECT 0.090 13.140 595.700 14.300 ;
        RECT 0.090 10.940 598.550 13.140 ;
        RECT 0.090 9.780 0.700 10.940 ;
        RECT 4.300 9.780 598.550 10.940 ;
        RECT 0.090 7.580 598.550 9.780 ;
        RECT 0.090 6.420 595.700 7.580 ;
        RECT 0.090 4.220 598.550 6.420 ;
        RECT 0.090 3.060 0.700 4.220 ;
        RECT 4.300 3.060 598.550 4.220 ;
        RECT 0.090 0.860 598.550 3.060 ;
        RECT 0.090 0.140 595.700 0.860 ;
      LAYER Metal4 ;
        RECT 36.540 21.930 98.740 571.670 ;
        RECT 100.940 21.930 175.540 571.670 ;
        RECT 177.740 21.930 252.340 571.670 ;
        RECT 254.540 21.930 329.140 571.670 ;
        RECT 331.340 21.930 405.940 571.670 ;
        RECT 408.140 21.930 482.740 571.670 ;
        RECT 484.940 21.930 559.540 571.670 ;
        RECT 561.740 21.930 588.420 571.670 ;
  END
END tiny_user_project
END LIBRARY

