* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_100_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5968__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout56_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _0012_ net80 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4640__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _0346_ net189 mod.pc0\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6776_ _0280_ net126 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3988_ _0951_ _0954_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_22_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5727_ mod.registers.r9\[5\] _2542_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _2442_ _2492_ _2497_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4609_ _0948_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5589_ _2403_ _2453_ _2455_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3903__B1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5504__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6629__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3682__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4564__B _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4698__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__B _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__B2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _3153_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4622__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ mod.registers.r3\[4\] _3165_ _0697_ mod.registers.r1\[4\] _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4891_ mod.instr_2\[5\] _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6630_ _0134_ net128 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5178__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3842_ _0801_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6561_ mod.des.des_dout\[18\] net3 _3124_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3773_ _0518_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5512_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ mod.des.des_dout\[7\] net5 _3080_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4138__B1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5443_ _2331_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ mod.registers.r2\[2\] _2304_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4325_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout105 net108 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout116 net119 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout127 net133 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout138 net143 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _0773_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ mod.registers.r1\[10\] _0697_ _0980_ mod.registers.r13\[10\] _1157_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6921__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _0332_ net122 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _0263_ net105 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A3 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4559__B _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3352__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3352__B2 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__I0 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3407__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4604__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4907__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5580__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout106_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ mod.registers.r3\[5\] _0471_ _0466_ mod.registers.r1\[5\] _3201_ mod.registers.r11\[5\]
+ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_96_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5090_ mod.pc0\[8\] _1892_ _1901_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4041_ _3215_ _3168_ mod.registers.r8\[7\] _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4943_ _1787_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ _1807_ _1832_ _1113_ _0711_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6613_ _0117_ net131 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3825_ mod.registers.r9\[15\] _0751_ _0730_ mod.registers.r10\[15\] _0795_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ mod.registers.r15\[14\] _3113_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3756_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5571__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ mod.des.des_counter\[0\] mod.des.des_counter\[1\] mod.des.des_counter\[2\]
+ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3687_ mod.registers.r5\[3\] _0547_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5426_ mod.registers.r3\[5\] _2338_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6520__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4126__A3 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5357_ _0958_ _2224_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3885__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0840_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ mod.pc_2\[7\] _2221_ _2224_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4239_ mod.registers.r4\[12\] _0971_ _0972_ mod.registers.r10\[12\] _1209_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3302__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4561__C _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6817__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__I _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3573__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3573__B2 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6511__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A2 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6967__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3628__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A1 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3610_ mod.pc_2\[5\] _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4590_ _1308_ _1311_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3541_ _0427_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6260_ mod.des.des_dout\[12\] _2921_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3472_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5305__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3316__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5211_ _2150_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6191_ _2857_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3867__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ _1924_ _2091_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5073_ _2032_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ mod.registers.r14\[14\] _0977_ _0978_ mod.registers.r7\[14\] _0981_ mod.registers.r9\[14\]
+ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4292__A2 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ mod.registers.r14\[14\] _2701_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _1824_ _1806_ _0661_ _1825_ _0429_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_138_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6592__I1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _1720_ _1727_ _1737_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_107_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _2413_ _3100_ _3105_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4888__I _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3739_ mod.registers.r14\[3\] _0607_ _0608_ mod.registers.r13\[3\] _0708_ _0709_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_119_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6458_ _2716_ _3062_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5409_ _2150_ _2327_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6389_ _2075_ _3009_ _3015_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__I _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5480__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6343__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6583__I1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__B2 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A1 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__B _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6518__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4274__A2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout173_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__B1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _2295_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3785__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _1098_ _1100_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3785__B2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5691_ _2425_ _2515_ _2519_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _0900_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4329__A3 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6574__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3537__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3537__B2 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4573_ _1531_ _1536_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2961_ _2965_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3524_ _3254_ _0470_ _0488_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ mod.instr\[8\] _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3455_ mod.instr_2\[11\] _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _1944_ _2859_ _2865_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout86_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3386_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ mod.pc\[10\] _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6428__I _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _2016_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5462__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _0607_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3473__B1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3787__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _2413_ _2688_ _2693_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _1826_ _1822_ _1824_ _1825_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5889_ mod.registers.r12\[14\] _2647_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3528__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3700__A1 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3700__B2 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__C _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__I0 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A1 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5756__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6181__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5444__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6492__I0 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6930_ _0028_ net164 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _0362_ net181 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5812_ _2527_ _2599_ _2602_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6792_ _0296_ net107 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3400__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5747__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _2260_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _2501_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4625_ _1350_ _1591_ _1593_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4183__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4183__B2 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _0593_ _1353_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ _3181_ _3162_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _1128_ _1151_ _1274_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _2899_ _2901_ _2902_ _2892_ _2898_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3438_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5683__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4486__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2851_ _2132_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _3192_ _3200_ _3205_ _3221_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5062__I _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3694__B1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ _2041_ _2065_ _2068_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6088_ _1959_ _2790_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5435__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4238__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5039_ _1989_ _2003_ net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4410__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5910__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput20 net20 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput31 net31 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4477__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_223 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_234 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_245 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_256 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5426__A1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_267 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_278 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_289 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5977__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3988__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4316__I _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout136_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4410_ _0992_ _1377_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ mod.registers.r2\[8\] _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4341_ _0757_ _0861_ _0650_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _2723_ mod.pc0\[1\] _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4468__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3676__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__C1 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__A1 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _0011_ net80 mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout49_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ _0345_ net181 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6393__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ _0279_ net104 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3987_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5726_ _2217_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3600__B1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ mod.registers.r7\[15\] _2493_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6850__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4156__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _3250_ _1558_ _1571_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5588_ mod.registers.r6\[4\] _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3903__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3903__B2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ _0918_ _1505_ _1508_ _1149_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3305__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6081__A1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4136__I _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4631__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6552__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3975__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__B _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6384__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4698__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5647__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4474__C _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6072__A1 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6723__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4622__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3425__A3 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3910_ mod.registers.r7\[4\] _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4890_ _1855_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ _0622_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6261__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _3125_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3772_ mod.registers.r5\[12\] _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _2193_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6491_ _3083_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__A2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4138__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4138__B2 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _2329_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5886__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ _2186_ _2302_ _2306_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _1288_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout106 net108 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout117 net119 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5638__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout128 net132 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout139 net143 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _1184_ _1190_ _1204_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4186_ _1153_ _1154_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6436__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__A2 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__B1 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _0331_ net122 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3795__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ _0262_ net101 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6689_ _0193_ net47 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__A1 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5515__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__A4 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3888__B1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3352__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4301__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4152__I1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__B1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5801__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6896__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4907__A3 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4540__A1 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5096__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ _0476_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2706_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1389_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6205__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _1826_ _1834_ _1835_ _1822_ _1825_ _1832_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_60_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6612_ _0116_ net76 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3824_ mod.registers.r1\[15\] _0746_ _0431_ mod.registers.r3\[15\] _0794_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5020__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6543_ _2435_ _3112_ _3115_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3755_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3686_ _0652_ _0653_ _0654_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6474_ _3072_ _3073_ _2789_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2205_ _2337_ _2339_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5356_ _2168_ _2107_ _1377_ _2273_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_114_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6769__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _1161_ _1164_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _2181_ _2024_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__A2 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _1136_ _1206_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4395__B _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ mod.registers.r3\[8\] _1013_ _1015_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6036__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4414__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3573__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5245__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5078__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__B1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3368__C _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5002__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout216_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ _0501_ _0504_ _0507_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4761__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3471_ _0415_ _0416_ _3289_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _2155_ _2157_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3316__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ _2867_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__I _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5141_ _2092_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5072_ mod.pc0\[7\] _1960_ _1961_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4023_ mod.registers.r4\[14\] _0971_ _0975_ mod.registers.r1\[14\] _0972_ mod.registers.r10\[14\]
+ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_111_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3403__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6018__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _2435_ _2700_ _2703_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5241__A2 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4925_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4234__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4856_ mod.ldr_hzd\[7\] _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3807_ _0498_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4787_ _1743_ _1747_ _1748_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6526_ mod.registers.r15\[7\] _3101_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4752__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3738_ _0660_ _3213_ _3214_ _3218_ _0662_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_118_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6457_ _1810_ _3058_ _3059_ _3041_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3669_ _0424_ _0636_ mod.registers.r4\[2\] _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5408_ _2160_ _2298_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6388_ mod.pc_1\[10\] _3010_ _3012_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ mod.registers.r1\[12\] _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _0107_ net209 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3313__I _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__B _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3794__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6934__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6248__A1 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3482__B2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout166_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _1678_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3785__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4982__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5690_ mod.registers.r8\[10\] _2516_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ _0878_ _1341_ _0716_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3537__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _0900_ _1537_ _1540_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6311_ mod.instr_2\[4\] _2958_ _2963_ mod.instr\[4\] _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3523_ _0489_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3454_ _3267_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6242_ _2912_ _2913_ _2914_ _2905_ _2911_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ mod.pc_1\[2\] _2861_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3385_ _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4657__C _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ _1914_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout79_I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ mod.pc0\[6\] _1960_ _1961_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6807__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ mod.registers.r11\[15\] _0974_ _0975_ mod.registers.r1\[15\] _0976_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5462__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3473__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3473__B2 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ mod.registers.r14\[7\] _2689_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1820_ _1819_ _1818_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5888_ _2564_ _2646_ _2649_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4839_ _1808_ _0445_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3528__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6509_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4489__B1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5150__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5453__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4110__C1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__I1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3464__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4716__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__C1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5692__A2 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5444__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6492__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _0361_ net193 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5811_ mod.registers.r11\[0\] _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6791_ _0295_ net107 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4404__B1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5742_ _2554_ _2551_ _2555_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _2400_ _2502_ _2508_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4707__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4624_ _0691_ _0808_ _0790_ _0800_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_135_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3915__C1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _0529_ _0681_ _0839_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3506_ _3175_ _3217_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3930__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4486_ _1448_ _1453_ _1454_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5132__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ mod.des.des_dout\[3\] _2896_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3437_ _3267_ _3269_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5683__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6156_ _2130_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3368_ mod.registers.r14\[0\] _3208_ _3211_ mod.registers.r13\[0\] _3220_ _3221_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_58_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__B2 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5107_ _2066_ _1891_ _2067_ _2041_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ _2782_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3299_ _0000_ mod.des.des_counter\[1\] _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6483__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _3223_ _1990_ _2002_ _1904_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input11_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5199__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _0087_ net221 mod.des.des_dout\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3749__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6123__B _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4174__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3685__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_224 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_235 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_246 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_257 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_268 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_279 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4332__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout129_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6652__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ _1059_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6259__I mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4271_ _0908_ _0910_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _2140_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__B2 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4873__C2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6912_ _0010_ net80 mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6843_ _0344_ net188 mod.pc0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__A1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _0278_ net103 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _0955_ _0952_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5725_ _2540_ _2541_ _2543_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3600__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5338__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3600__B2 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5656_ _2439_ _2492_ _2496_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _1572_ _1556_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5587_ _2447_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3903__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4538_ _1506_ _0934_ _1507_ _1484_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__B1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4469_ _1337_ _1251_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6208_ _2717_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6139_ _2828_ _2827_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6118__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__A1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A1 _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3940__B _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A3 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3830__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ _0776_ _0803_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _0517_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5510_ _2394_ _2389_ _2395_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6490_ mod.des.des_dout\[6\] net4 _3080_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5441_ _2268_ _2343_ _2348_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5335__A1 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5886__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5372_ mod.registers.r2\[1\] _2304_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4323_ _1203_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5638__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout129 net132 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4254_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4438__S _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4310__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ mod.registers.r12\[10\] _1110_ _1106_ mod.registers.r10\[10\] _1155_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4861__A3 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5271__B1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__B2 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _0330_ net105 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _0261_ net106 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3969_ _3233_ _0926_ _3249_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _2528_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6688_ _0192_ net90 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__A1 _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _2472_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5877__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3888__B2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6054__A2 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6563__S _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__B2 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__B2 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4907__A4 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3576__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A1 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3654__C _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3879__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout196_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6840__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5990_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4056__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _1909_ _1578_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4851__I0 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _1824_ _1836_ _0616_ _0951_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6611_ _0115_ net77 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6990__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ mod.registers.r6\[15\] _0733_ _0766_ mod.registers.r12\[15\] _0793_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3406__I1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3567__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ mod.registers.r15\[13\] _3113_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3754_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _2966_ _3044_ _3066_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3685_ mod.registers.r4\[3\] _0508_ _0421_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5424_ mod.registers.r3\[4\] _2338_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _2270_ _2290_ _2291_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4306_ _1259_ _1271_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5286_ _2201_ _2229_ _2230_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4237_ _0956_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4295__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4168_ mod.registers.r15\[8\] _0963_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4047__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4099_ _1067_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5244__B1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3739__C _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6809_ _0313_ net118 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4430__I _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6713__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4286__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__B2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6027__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3797__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3549__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4340__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3470_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout209_I net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5710__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3316__A3 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _2094_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A3 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6267__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5071_ _2033_ _1963_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4029__B2 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ mod.registers.r14\[13\] _2701_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4515__I _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _1388_ _1787_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4855_ mod.ldr_hzd\[4\] _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3806_ _0756_ _0775_ _0496_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _1749_ _1753_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6736__CLK net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _2410_ _3100_ _3104_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3737_ mod.registers.r11\[3\] _0705_ _0706_ mod.registers.r8\[3\] _0707_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5346__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _2992_ _3061_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3668_ _0637_ _0633_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5407_ _2296_ _2321_ _2326_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5701__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4504__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _0862_ _3009_ _3014_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6886__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3599_ mod.registers.r4\[4\] _0420_ _0449_ mod.registers.r1\[4\] _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5338_ _2178_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6257__A2 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _1078_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ _0106_ net209 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4853__C _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5768__A1 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3779__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__I0 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6193__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A4 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6248__A2 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3482__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4335__I _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout159_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _0809_ _0842_ _0876_ _0725_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _1241_ _1338_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__I _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _2961_ _2964_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3522_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6241_ mod.des.des_dout\[7\] _2909_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3453_ _3280_ _3288_ _0414_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_103_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ _2753_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3384_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5123_ _2056_ _2074_ _2080_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _2017_ _1963_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4005_ _3178_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3473__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4670__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5956_ _2410_ _2688_ _2692_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4907_ _1802_ _1810_ _1804_ _1807_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5887_ mod.registers.r12\[13\] _2647_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4973__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__A1 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _0637_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5922__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _1280_ _1652_ _1651_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _3091_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _3048_ _3049_ _3046_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4489__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__B2 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5150__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__B1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__C2 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3464__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6901__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6402__A2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__I _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6370__I _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5913__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__B1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__C2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4774__B _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5810_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6790_ _0294_ net103 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4404__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4404__B2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5741_ mod.registers.r9\[9\] _2552_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ mod.registers.r8\[3\] _2504_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6213__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _1409_ _1592_ _1344_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5904__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3409__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3915__B1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3915__C2 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4554_ _1344_ _1356_ _1364_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_156_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5380__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3505_ mod.registers.r11\[1\] _3202_ _3195_ mod.registers.r10\[1\] _0475_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4485_ _1097_ _1049_ _1249_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout91_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5132__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ mod.instr_2\[11\] _3276_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6155_ _2833_ _2838_ _2841_ _2847_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ _3212_ _3213_ _3214_ _3218_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_98_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3694__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5106_ mod.pc0\[9\] _1891_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1943_ _2784_ _1959_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4684__B _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3298_ mod.des.des_counter\[0\] _3150_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6924__CLK net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _1998_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4643__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5199__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6396__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6988_ _0086_ net216 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5939_ _2679_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3749__A3 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6148__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4159__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4174__A3 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3382__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5534__I _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5123__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3685__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3989__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_225 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_236 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_247 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_258 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_269 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6387__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5709__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__B1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4270_ _1004_ _1238_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6311__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__B2 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6947__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4873__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4873__B2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6275__I mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4625__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _0009_ net81 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6842_ _0343_ net186 mod.pc0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3848__B _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ _0277_ net126 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ mod.funct7\[2\] _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5050__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5724_ mod.registers.r9\[4\] _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3600__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5655_ mod.registers.r7\[14\] _2493_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4606_ _1366_ _1573_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ _2445_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4537_ _1506_ _1349_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__C _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6302__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _1253_ _1099_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6302__B2 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6207_ mod.instr\[0\] _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3419_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4399_ _0934_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6138_ _1913_ _2083_ _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _1926_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4616__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5529__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6541__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4147__A3 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4589__B _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3940__C _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3512__I _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5280__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout141_I net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3770_ _0731_ _0734_ _0737_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5583__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ mod.registers.r3\[11\] _2344_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6532__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5371_ _2177_ _2302_ _2305_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _1291_ _1220_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5099__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout119 net123 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4253_ _1221_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3649__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ mod.registers.r5\[10\] _0882_ _0696_ mod.registers.r4\[10\] _0706_ mod.registers.r8\[10\]
+ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4310__A3 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout54_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5271__A1 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3821__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _0329_ net119 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5023__A1 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6756_ _0260_ net70 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3968_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3585__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5707_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6687_ _0191_ net53 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3899_ mod.registers.r13\[9\] _0541_ _0542_ mod.registers.r1\[9\] _0869_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6523__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _2414_ _2480_ _2485_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5569_ _2295_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3576__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3576__B2 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3879__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4828__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout189_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5253__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _3243_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__I1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__B mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4871_ _1839_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3822_ mod.registers.r5\[15\] _0440_ _0442_ mod.registers.r7\[15\] _0792_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _0114_ net77 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3567__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _2430_ _3112_ _3114_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3567__B2 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3753_ _0719_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6505__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _1820_ _3064_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5308__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3684_ mod.registers.r11\[3\] _0505_ _0506_ mod.registers.r2\[3\] _0654_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6221__C _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _2331_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5354_ mod.registers.r1\[14\] _2277_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4305_ _1127_ _1150_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ mod.registers.r1\[6\] _2206_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4819__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ _1044_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5492__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6665__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4167_ _1135_ _1136_ mod.registers.r1\[8\] _1015_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ _0759_ _0494_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4047__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__B2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _0312_ net101 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6739_ _0243_ net69 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__C _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4286__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6574__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3997__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5235__A1 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__B2 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3549__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3549__B2 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout90 net94 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4210__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout104_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5452__I _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ mod.pc\[7\] _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5474__A1 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ _0988_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _2430_ _2700_ _2702_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6216__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4923_ mod.pc\[0\] _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4017__B _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ mod.ldr_hzd\[5\] _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ _0757_ _0773_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4785_ _1167_ _1669_ _1754_ _1659_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4531__I _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ mod.registers.r15\[6\] _3101_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3736_ _3204_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3667_ _0425_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6455_ _1804_ _3058_ _3059_ _3036_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ mod.registers.r2\[15\] _2322_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6386_ mod.pc_1\[9\] _3010_ _3012_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4687__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3598_ mod.registers.r10\[4\] _3279_ _0413_ mod.registers.r2\[4\] _0568_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3712__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5337_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5268_ _2172_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6501__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7007_ _0105_ net210 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4219_ _1185_ _1188_ _1181_ _1165_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _2146_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6407__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3610__I mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4440__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6568__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6142__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__I _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3951__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6830__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3703__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__I _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4259__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6980__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5208__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3520__I mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout221_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4195__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _0989_ _1538_ _1422_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5931__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _0490_ _0482_ _3258_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6479__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _2718_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ mod.registers.r4\[0\] _0420_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6171_ _2781_ _2859_ _2863_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3383_ _3234_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5122_ _2005_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5447__A1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ mod.pc\[6\] _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4004_ _0605_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3430__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5955_ mod.registers.r14\[6\] _2689_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _1831_ _1847_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5886_ _2560_ _2646_ _2648_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ mod.ldr_hzd\[8\] _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4261__I _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _1281_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5922__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3719_ _0470_ _0488_ _0560_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4699_ _0945_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _2967_ _1862_ _3038_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__A1 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__B _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6369_ _0651_ _3000_ _3002_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5438__A1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__A1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4110__B2 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6137__B mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3621__B1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4177__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A2 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3924__B2 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5677__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6047__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout171_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3860__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5601__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _2253_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6876__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3612__B1 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5671_ _2397_ _2502_ _2507_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4168__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4622_ _0529_ _0773_ _0681_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_135_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3915__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3915__B2 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4553_ _1383_ _1513_ _1516_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_156_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3504_ mod.registers.r8\[1\] _0473_ _3199_ mod.registers.r9\[1\] _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4484_ _1269_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5668__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _2717_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3435_ mod.registers.r14\[0\] _3283_ _3287_ mod.registers.r6\[0\] _3288_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ _2774_ _2848_ _2849_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3366_ mod.registers.r15\[0\] _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout84_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5105_ mod.pc\[9\] _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6085_ _2768_ _2769_ mod.pc\[3\] _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3297_ _3152_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5640__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5036_ mod.pc0\[5\] _1960_ _1961_ _2000_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_73_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4643__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4256__I _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _0085_ net216 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6396__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5938_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6404__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5869_ mod.registers.r12\[6\] _2635_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4159__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4159__B2 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3906__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3382__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput23 net23 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_226 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6084__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_237 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_248 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_259 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5831__A1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__I _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4398__B2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5898__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4570__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _0008_ net81 mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6492__S _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6841_ _0342_ net180 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4389__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _0276_ net71 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3984_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5723_ _2531_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ _2436_ _2492_ _2495_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5889__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _1555_ _1349_ _1371_ _1450_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5585_ _2400_ _2446_ _2452_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4561__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ _1148_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _1097_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6206_ _2131_ _2883_ _2886_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4313__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3418_ _3267_ _3269_ _3270_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4398_ _1362_ _1363_ _1365_ _0627_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _2802_ _1885_ mod.pc\[10\] _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3349_ _3201_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _1911_ _2004_ _1920_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4077__B1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4616__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ _3153_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A3 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6415__B _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6541__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__I _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__B1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5804__A1 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__B1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3949__B _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4240__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6532__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ mod.registers.r2\[0\] _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4321_ mod.pc_2\[12\] _1205_ _1289_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5099__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4252_ _0755_ _1220_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_86_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4183_ mod.registers.r15\[10\] _0884_ _0879_ mod.registers.r7\[10\] mod.registers.r3\[10\]
+ _0694_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_80_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5190__I _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4059__B1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__C _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5271__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout47_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _0328_ net97 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ _0259_ net70 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3967_ _0931_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5706_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3585__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4782__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6686_ _0190_ net48 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3898_ mod.registers.r15\[9\] _0435_ _0437_ mod.registers.r12\[9\] _0868_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5637_ mod.registers.r7\[7\] _2481_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4534__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ _2439_ _2432_ _2440_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4519_ _1462_ _1465_ _1466_ _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5499_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6287__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3648__I0 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__C _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__B _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3576__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6514__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6278__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4828__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A2 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__I2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4870_ _1815_ _1834_ _1836_ _1813_ _1812_ _1832_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_3821_ mod.registers.r13\[15\] _0745_ _0732_ mod.registers.r14\[15\] _0791_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6540_ mod.registers.r15\[12\] _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3567__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4764__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3752_ _3239_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _3070_ _3071_ _3057_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6505__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3683_ mod.registers.r14\[3\] _0534_ _0535_ mod.registers.r6\[3\] _0653_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5422_ _2329_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4516__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4304_ _1272_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5284_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4819__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4235_ _0778_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5492__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _0483_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ mod.pc_2\[1\] _0777_ _1065_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4047__A3 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6441__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _0311_ net106 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4055__I0 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1959_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _0242_ net69 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _0173_ net52 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5095__I _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3608__I _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4507__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3343__I _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3549__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net81 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net94 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4123__B _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5474__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _0989_ _0986_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3485__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__B _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ mod.registers.r14\[12\] _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4985__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _1822_ _1809_ _0636_ _0424_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4737__A1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__C1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ _0552_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4784_ _1400_ _1595_ _1481_ _1317_ _1660_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _2407_ _3100_ _3103_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3735_ _3202_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4033__B _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _2992_ _3060_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3666_ _0562_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5405_ _2290_ _2321_ _2325_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6385_ _0843_ _3009_ _3013_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3597_ _0558_ _0559_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6632__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3712__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5336_ mod.des.des_dout\[33\] _2248_ _2272_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_115_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _2165_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7006_ _0104_ net206 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4218_ _1186_ _1187_ _1126_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3476__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6782__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _2147_ _2143_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ mod.registers.r15\[9\] _0884_ _0600_ mod.registers.r6\[9\] _0473_ mod.registers.r8\[9\]
+ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4189__C1 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3338__I _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3951__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3703__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6585__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6405__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4118__B _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3957__B _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4195__A2 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3520_ mod.instr_2\[4\] _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3451_ _3236_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ mod.pc_1\[1\] _2861_ _2822_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3382_ _3230_ _3231_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4079__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5121_ _2060_ _2078_ _2076_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_151_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6495__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5447__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ _1911_ _2004_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5998__A3 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6294__I _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4003_ mod.registers.r4\[15\] _0971_ _0972_ mod.registers.r10\[15\] _0973_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3711__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4958__B2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _2407_ _2688_ _2691_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4970__C _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4905_ _1831_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5885_ mod.registers.r12\[12\] _2647_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4836_ _3275_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5383__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _1728_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3718_ _0687_ _0492_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _1665_ _1666_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6437_ _1825_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3649_ _0615_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5686__A2 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6368_ mod.pc_1\[3\] _3001_ _2996_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3697__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4894__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4894__C2 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ mod.des.des_dout\[31\] _2248_ _2257_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6299_ _0905_ _2956_ _2951_ mod.instr\[0\] _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6486__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4949__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__B _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3621__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5548__I _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3621__B2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5374__A1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4177__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5677__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3688__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4101__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3860__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3860__B2 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout164_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3612__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__I _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3612__B2 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4362__I _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ mod.registers.r8\[2\] _2504_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4168__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _0827_ _0841_ _0802_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3915__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4552_ _1520_ _1521_ _1432_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _3203_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4483_ _1449_ _1451_ _1452_ _1445_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5193__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5668__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ mod.instr\[3\] _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3434_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6153_ mod.pc\[12\] _2774_ _2822_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3365_ _3215_ _3216_ _3209_ _3217_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_98_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _2056_ _2055_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _1944_ _2780_ _2787_ _2789_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3296_ net176 _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6093__A2 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _1999_ _1963_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4643__A3 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3851__A1 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3851__B2 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6986_ _0084_ net216 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6820__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__I _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3603__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4272__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _2544_ _2634_ _2637_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6970__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4159__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _0902_ _1785_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5799_ _2560_ _2591_ _2593_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3367__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3906__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4867__C2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_227 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_238 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6084__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_249 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5595__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4182__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3526__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4322__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ _0341_ net180 mod.pc0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6993__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6771_ _0275_ net74 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3983_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5722_ _2529_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ mod.registers.r7\[13\] _2493_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5916__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__I _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _1068_ _0933_ _0939_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5584_ mod.registers.r6\[3\] _2448_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ _1327_ _0810_ _0877_ _1339_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4561__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4466_ _1242_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ mod.pc_1\[13\] _2884_ _2880_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5510__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ mod.instr_2\[11\] mod.instr_2\[10\] _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4313__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _2833_ _2829_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3348_ _3196_ _3197_ _3160_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4077__B2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5018_ _1969_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3824__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _0067_ net217 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3588__B1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5329__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6716__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3346__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__B2 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5568__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3579__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4240__B2 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4791__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout127_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _0742_ _0744_ _0750_ _0753_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_153_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3897__A4 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4796__B _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__I _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4251_ _0755_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4182_ _0489_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6048__A2 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4059__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4059__B2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _0327_ net98 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5559__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _0258_ net70 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4231__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3966_ _3226_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4231__B2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _2161_ _2499_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ _0189_ net52 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4782__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _0863_ _0864_ _0865_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_136_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ _2411_ _2480_ _2484_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5567_ mod.registers.r5\[14\] _2433_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5731__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ _1224_ _1397_ _1479_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _2176_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4449_ _0715_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4298__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6119_ _2033_ _2780_ _2819_ _2789_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5798__A1 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3648__I1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6426__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6598__I0 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4222__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__B2 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__I _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5789__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__I3 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ _0779_ _0789_ _0556_ _0557_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_33_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3751_ _0720_ _0712_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5961__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4764__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _3055_ _3041_ _3066_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3682_ mod.registers.r8\[3\] _0531_ _0532_ mod.registers.r10\[3\] _0652_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _2199_ _2330_ _2336_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5713__A1 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4516__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5352_ mod.des.des_dout\[35\] _2220_ _2286_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_99_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ _1180_ _1181_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6297__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5283_ mod.des.des_dout\[27\] _2220_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3714__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _3183_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _0675_ _0676_ _0677_ _0678_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4452__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _0310_ net101 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4204__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ mod.pc0\[3\] _1960_ _1961_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4055__I1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6737_ _0241_ net45 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5952__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ _0718_ _0913_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _0172_ net142 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ _2471_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6599_ _3147_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6904__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout70 net72 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout81 net82 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout92 net94 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_127_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3706__B1 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5235__B _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__A1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout194_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3485__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _2682_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4985__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6580__I _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6187__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ mod.ldr_hzd\[6\] _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4198__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3803_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4198__C2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4737__A2 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _1750_ _1751_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6522_ mod.registers.r15\[5\] _3101_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ mod.registers.r10\[3\] _0602_ _0703_ mod.registers.r9\[3\] _0704_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _1807_ _3058_ _3059_ _1862_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3665_ _0631_ _0632_ mod.registers.r11\[2\] _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ mod.registers.r2\[14\] _2322_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6384_ mod.pc_1\[8\] _3010_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3596_ mod.registers.r13\[4\] _0447_ _0431_ mod.registers.r3\[4\] _0565_ _0566_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_161_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5335_ _2025_ _2273_ _2166_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3712__A3 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6111__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _0580_ _2189_ _2209_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6927__CLK net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7005_ _0103_ net206 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4217_ _0859_ _1147_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5197_ mod.rd_3\[3\] _2144_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3476__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4673__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _1114_ _1115_ _1116_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6414__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4079_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3779__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5925__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__C2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4900__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4113__B1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6405__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3529__I _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4195__A3 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3450_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout207_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3381_ mod.instr_2\[1\] _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _2077_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ _2005_ _2007_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4655__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4002_ _0602_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ mod.registers.r14\[5\] _2689_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _1866_ _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5884_ _2628_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4835_ _0633_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3439__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5383__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _1332_ _1731_ _1732_ _1735_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6505_ _2327_ _2624_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3717_ _0615_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4697_ _1307_ _1544_ _0922_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _3032_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3648_ mod.instr_2\[5\] _0616_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6367_ _2952_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3579_ mod.registers.r5\[7\] _0547_ _0548_ mod.registers.r7\[7\] _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3697__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4894__B2 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ _2174_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6298_ _2955_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6485__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _0651_ _2168_ _2173_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4646__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4219__B _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4949__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5071__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5829__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3349__I _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5374__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3793__B _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3688__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4637__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3860__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6622__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout157_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3612__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4620_ _1267_ _1349_ _0921_ _1587_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5365__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1438_ _1519_ _1495_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3502_ mod.registers.r3\[1\] _0471_ _3186_ mod.registers.r6\[1\] mod.registers.r7\[1\]
+ _3170_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_143_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4482_ _1056_ _1061_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _2895_ _2719_ _2897_ _2892_ _2898_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3433_ _3284_ _3285_ _3274_ _3276_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6152_ _2845_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _3159_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _2059_ _2062_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6083_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3295_ _0000_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6238__C _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ mod.pc\[5\] _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3300__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3851__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _0083_ net116 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5649__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _2299_ _2624_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3603__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ mod.registers.r12\[5\] _2635_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4818_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5356__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ mod.registers.r10\[12\] _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3906__A3 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4749_ _1713_ _1714_ _1715_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_119_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5108__A2 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _1812_ _0003_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xoutput25 net25 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput36 net36 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4867__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4867__B2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5333__B _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3632__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_228 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_239 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3827__C1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4095__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__A4 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4463__I _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6795__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5347__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3807__I _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3542__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__A1 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__S _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6770_ _0274_ net71 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3982_ _3232_ _3252_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _2204_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6535__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _2431_ _2492_ _2494_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4603_ _1309_ _1333_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5583_ _2397_ _2446_ _2451_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4534_ _1420_ _1502_ _1503_ _0920_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6299__B1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4465_ _1398_ _1428_ _1431_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_104_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _2115_ _2883_ _2885_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3416_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4396_ _0725_ _0920_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6135_ _2816_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4548__I _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3347_ mod.registers.r10\[0\] _3195_ _3199_ mod.registers.r9\[0\] _3200_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6668__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _2726_ _1900_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5017_ _1979_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4283__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6968_ _0066_ net217 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3588__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3588__B2 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5919_ _2416_ _2667_ _2669_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4785__B1 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6899_ _0400_ net164 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6526__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6129__I1 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6159__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3362__I _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4068__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5017__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3579__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__B2 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4240__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4250_ _1205_ _1208_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6960__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5008__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6822_ _0326_ net93 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5559__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _0257_ net69 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5927__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ mod.funct3\[0\] _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3648__S _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4231__A2 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _2176_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6684_ _0188_ net114 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3896_ mod.registers.r4\[9\] _0508_ _0421_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5635_ mod.registers.r7\[6\] _2481_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5566_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5731__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4517_ _1332_ _1483_ _1486_ _1222_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5662__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5497_ _2296_ _2379_ _2384_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4448_ _1400_ _1408_ _1417_ _1329_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5495__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4379_ _3229_ _3244_ _3247_ _0936_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6118_ _2814_ _2817_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5247__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6049_ _2741_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6598__I1 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6442__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6161__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6833__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3497__B1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4461__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3976__B _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3750_ _0560_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ mod.pc_2\[3\] _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_158_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5420_ mod.registers.r3\[3\] _2332_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _2220_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4302_ _1165_ _1166_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5282_ _2222_ _2223_ _2225_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5477__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4233_ _0772_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _0711_ _1113_ mod.registers.r8\[8\] _1010_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5229__A1 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3730__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _0670_ _0671_ _0672_ _0673_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6246__C _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout52_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6706__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4452__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3660__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _0309_ net105 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _1962_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4204__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5401__A1 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6856__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0240_ net62 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3948_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4755__A3 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6667_ _0171_ net142 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3879_ mod.registers.r12\[8\] _0848_ _0638_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5618_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6598_ net6 mod.des.des_dout\[34\] _3136_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5549_ mod.registers.r5\[10\] _2419_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4691__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5943__A2 _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout71 net72 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3706__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__B2 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4131__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3485__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout187_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4920_ _1884_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6879__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3642__B1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _1817_ _1818_ _1819_ _1820_ _1805_ _1808_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6187__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4381__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3802_ _0758_ _0759_ _0764_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4198__B2 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4782_ _1467_ _1587_ _1329_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6521_ _2402_ _3100_ _3102_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3733_ _3198_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _2147_ _2966_ _3025_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3664_ _0444_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5698__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2284_ _2321_ _2324_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6383_ _2752_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3595_ _0560_ _0561_ _0563_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5334_ _2224_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6111__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ _2210_ _1988_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _0102_ net205 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4216_ _0874_ _1124_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5196_ _1848_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5870__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3476__A3 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4673__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4147_ _0951_ _0616_ mod.registers.r4\[9\] _1010_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4078_ _0524_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5622__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4505__B _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4189__B2 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _0223_ net54 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3635__I _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4113__A1 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4113__B2 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4466__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3370__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5613__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3545__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout102_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5760__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1790_ _2013_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4104__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5301__B1 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ _3174_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5604__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _2402_ _2688_ _2690_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ mod.instr_2\[6\] _1869_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _2626_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4834_ mod.ldr_hzd\[9\] _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _1204_ _1397_ _1546_ _1330_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6504_ _3090_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3716_ _0682_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _1322_ _1355_ _0497_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6435_ _3043_ _3045_ _3046_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4060__B _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3647_ _3258_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _2713_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3578_ _0441_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4894__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1991_ _2226_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _2856_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5248_ _2169_ _1950_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5843__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4646__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _2072_ _2120_ _2134_ _3156_ _2135_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__B _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4889__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4582__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4885__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__B1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6917__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4550_ _1438_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_156_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ _3164_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4481_ _1068_ _1450_ _0454_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6220_ _2788_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3432_ mod.instr_2\[12\] _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6151_ _2114_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3363_ _3162_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ _2059_ _2062_ _1790_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3294_ mod.des.des_counter\[1\] _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _2706_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__B1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4628__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _1934_ _1912_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3300__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _0082_ net116 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6254__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5935_ _2441_ _2673_ _2678_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4800__A2 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5866_ _2540_ _2634_ _2636_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _0908_ _1784_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5665__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _2573_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5356__A3 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3367__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4564__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _1716_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _1259_ _1271_ _1492_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6349_ _0711_ _2989_ _2986_ mod.instr\[17\] _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5816__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_229 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3827__B1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__C2 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4095__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6445__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__A1 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5575__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5283__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3981_ _3196_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5720_ _2538_ _2530_ _2539_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5651_ mod.registers.r7\[12\] _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6090__B _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6535__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _1382_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5582_ mod.registers.r6\[2\] _2448_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4533_ _0924_ _0927_ _0717_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6299__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__B2 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4464_ _1302_ _1296_ _1399_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_117_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6203_ mod.pc_1\[12\] _2884_ _2880_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3415_ mod.instr_2\[12\] _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3733__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4395_ _1226_ _1357_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6249__C _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6134_ mod.pc\[10\] _2824_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout82_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _1893_ _2766_ _2772_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ mod.pc0\[4\] _1922_ _1923_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _0065_ net219 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ mod.registers.r13\[8\] _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3588__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__B2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6898_ _0399_ net164 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ _2355_ _2498_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3908__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4537__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6612__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4225__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3579__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4423__B _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3751__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4180_ _1148_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6453__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__B2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__B mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6205__A1 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5008__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__C _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6821_ _0325_ net97 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6752_ _0256_ net57 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3964_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ _2442_ _2521_ _2526_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4231__A3 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6683_ _0187_ net114 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4333__B _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3895_ mod.registers.r11\[9\] _3292_ _0506_ mod.registers.r2\[9\] _0865_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5634_ _2408_ _2480_ _2483_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5148__C _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5565_ _2289_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6635__CLK net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4516_ _1228_ _1369_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ mod.registers.r4\[15\] _2380_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3463__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4447_ _1400_ _1412_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5495__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ _1332_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6117_ _2764_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ mod.instr_2\[15\] _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6444__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6048_ _2730_ _2105_ _2758_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3497__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3497__B2 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4213__A3 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3548__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6658__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout132_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3680_ _0628_ _0577_ _0643_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_71_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _1233_ _2273_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ _1263_ _1268_ _1269_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5281_ _2171_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4232_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ mod.registers.r6\[8\] _0700_ _0696_ mod.registers.r4\[8\] _0603_ mod.registers.r9\[8\]
+ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4094_ _1055_ _1061_ _1062_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4328__B _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout45_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3660__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5938__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__B2 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6804_ _0308_ net73 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ _1924_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6262__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5401__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6735_ _0239_ net63 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3947_ _3227_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3458__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _0170_ net140 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3878_ _0631_ _0562_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5165__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _3146_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5548_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4912__B2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6114__B1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _2361_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3921__I _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6417__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A3 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__I _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout61 net65 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout72 net75 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout83 net88 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout94 net100 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6950__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6105__B1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4927__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3831__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6408__A1 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3642__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__B _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3642__B2 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ mod.ldr_hzd\[15\] _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3801_ _0767_ _0768_ _0769_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4198__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5395__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _1352_ _1404_ _1473_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ mod.registers.r15\[4\] _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3732_ mod.registers.r6\[3\] _0700_ _0468_ mod.registers.r5\[3\] mod.registers.r2\[3\]
+ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _3032_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6589__I _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _3276_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5698__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ mod.registers.r2\[13\] _2322_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6382_ _0530_ _3009_ _3011_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3594_ mod.registers.r15\[4\] _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5333_ _2123_ _2189_ _2214_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _1793_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _0101_ net205 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4215_ _1166_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3741__I _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _2141_ _2143_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5870__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4146_ _0482_ _0483_ mod.registers.r13\[9\] _0478_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4077_ _1021_ _1043_ _1046_ _0458_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_83_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5622__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4505__C _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4189__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5386__A1 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6973__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1943_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6718_ _0222_ net49 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6649_ _0153_ net138 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__B1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3872__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5613__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4352__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3561__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4000_ _0961_ _0965_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ mod.registers.r14\[4\] _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6093__B mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6996__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4902_ _1870_ _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5882_ _2558_ _2640_ _2645_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _1802_ _0429_ _0632_ _0846_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4764_ _0922_ _1733_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ mod.des.des_dout\[12\] net10 _3074_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3715_ _0683_ _0684_ _0453_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3736__I _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _1315_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6434_ _2715_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5156__C _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3646_ _3216_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _0628_ _2714_ _2999_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3577_ _0439_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _2075_ _2189_ _2209_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2951_ _2954_ _2831_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5247_ _2164_ _2194_ _2195_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _3154_ _2122_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4129_ _1093_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7001__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5398__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4516__B _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5359__A1 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4031__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6719__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4582__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__CLK net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3381__I mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4098__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3845__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4940__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5257__B _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A1 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3556__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ _0467_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout212_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4480_ _0688_ _0689_ _1069_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3431_ mod.instr_2\[13\] _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6570__I0 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6150_ mod.pc\[12\] _1914_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _3181_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5101_ _2060_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6081_ _2765_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3293_ mod.des.des_counter\[0\] _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__B2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _1915_ _1988_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5038__B1 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _0081_ net116 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ mod.registers.r13\[15\] _2674_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ mod.registers.r12\[4\] _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4816_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _2571_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4747_ _1030_ _1669_ _1485_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _1280_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6417_ _2728_ _1801_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5513__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _0597_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput27 net27 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput38 net38 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6348_ _2860_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ mod.instr\[17\] _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__B2 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6017__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6241__A2 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5752__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6691__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4307__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__S _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout162_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3980_ _0779_ _0878_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ _2474_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ _1563_ _1567_ _1570_ _0918_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5581_ _2394_ _2446_ _2450_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4546__A2 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4532_ _1500_ _1470_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6299__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4463_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _2857_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3414_ mod.instr_2\[13\] _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _0529_ _1291_ _0553_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6133_ _2825_ _2830_ _2831_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3345_ _3196_ _3197_ _3175_ _3187_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__I _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6064_ _2767_ _2771_ _2754_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout75_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _1980_ _1897_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6265__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _0064_ net217 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _2655_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4785__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ _0398_ net177 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _2568_ _2618_ _2623_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4537__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _2540_ _2579_ _2581_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6501__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__B2 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5973__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5725__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4464__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _0324_ net39 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4216__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6751_ _0255_ net42 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5964__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _0930_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4767__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ mod.registers.r8\[15\] _2522_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6682_ _0186_ net96 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3894_ mod.registers.r14\[9\] _0534_ _0535_ mod.registers.r6\[9\] _0864_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5716__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ mod.registers.r7\[5\] _2481_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5564_ _2436_ _2432_ _2437_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _2290_ _2379_ _2383_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4446_ _1351_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _1328_ _1335_ _1340_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6116_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3328_ _3161_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _2729_ mod.pc0\[11\] _2754_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6444__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4455__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6949_ _0047_ net149 mod.ldr_hzd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4524__B _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__I _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__I _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3497__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4694__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5946__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__A4 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout125_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3564__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4300_ _1033_ _1048_ _1094_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6123__A1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ _1046_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _1135_ _1191_ _0561_ _0985_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_99_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ mod.registers.r10\[8\] _1106_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6096__B _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ _0719_ _0722_ _0666_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_110_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6803_ _0307_ net73 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ mod.pc\[3\] _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6734_ _0238_ net58 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3946_ _0914_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6665_ _0169_ net140 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3877_ _0846_ _0632_ mod.registers.r11\[8\] _0634_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_109_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _2327_ _2356_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5165__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ net5 mod.des.des_dout\[33\] _3142_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6752__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _2260_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5478_ _2359_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4429_ _1237_ _1287_ _1295_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout40 net46 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout51 net56 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4600__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout62 net64 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout73 net75 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout84 net86 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5864__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout95 net99 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3384__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4116__B1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4667__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6408__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4943__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3642__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3559__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ mod.registers.r5\[13\] _0741_ _0743_ mod.registers.r7\[13\] _0770_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4780_ _1665_ _1415_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__CLK net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3731_ _3190_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3945__A3 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3662_ _0416_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5147__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6344__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _3054_ _3056_ _3057_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6344__B2 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ _2276_ _2321_ _2323_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6381_ mod.pc_1\[7\] _3010_ _3004_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3593_ _0415_ _0562_ _0444_ _3277_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_115_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _2210_ _2108_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5263_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7002_ _0100_ net205 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4214_ _1102_ _1105_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5194_ mod.rd_3\[2\] _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4145_ _0480_ _3256_ mod.registers.r14\[9\] _0478_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_28_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5014__I mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _1044_ _0491_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5386__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ mod.pc0\[2\] _1922_ _1923_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3397__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6717_ _0221_ net55 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5684__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3929_ _0759_ _0896_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_109_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _0152_ net127 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6335__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6335__B2 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3932__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__B2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__I0 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4821__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3624__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6798__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5301__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout192_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _2682_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3615__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4901_ mod.ldr_hzd\[8\] _1856_ _1858_ mod.ldr_hzd\[10\] mod.instr_2\[5\] _1871_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5881_ mod.registers.r12\[11\] _2641_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ mod.ldr_hzd\[11\] _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3379__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _1333_ _1365_ _0627_ _1359_ _1666_ _1343_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6502_ _3089_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3714_ _0557_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6317__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4694_ _1659_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _3029_ _3044_ _3038_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3645_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6364_ mod.pc_1\[2\] _2995_ _2996_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3576_ mod.registers.r9\[7\] _0544_ _0545_ mod.registers.r3\[7\] _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5315_ _2210_ _2074_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6295_ _1886_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ mod.registers.r1\[2\] _2179_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _2130_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _1076_ _1093_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5056__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ mod.pc_2\[7\] _0499_ _1027_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4803__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5359__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3790__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A1 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__CLK net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3430_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6570__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3361_ _3206_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ mod.pc_2\[9\] _1233_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6080_ _2783_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6963__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _1916_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _0080_ net116 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5589__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _2438_ _2673_ _2677_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5864_ _2628_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _0904_ _0905_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5795_ _2558_ _2585_ _2590_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _1031_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5761__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3772__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4677_ _1511_ _1554_ _1579_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6416_ _2147_ _2956_ _3031_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3628_ mod.registers.r4\[2\] _3174_ _3178_ mod.registers.r1\[2\] _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6561__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput28 net28 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6347_ _2985_ _2988_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3559_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _2939_ _2937_ _2940_ _2941_ _2935_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5277__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ mod.registers.r1\[0\] _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3827__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4252__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6836__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5752__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__A3 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6552__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6986__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3515__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3392__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6208__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__C1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__B1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5440__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout155_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _0726_ _1568_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5580_ mod.registers.r6\[1\] _2448_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4546__A3 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _1305_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4462_ _3250_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6201_ _2867_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3506__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3413_ _3265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4393_ _0925_ _1334_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6132_ _2707_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3344_ mod.instr_2\[16\] _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _1797_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ mod.pc\[4\] _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6709__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout68_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4482__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _0063_ net219 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5431__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _2653_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _0397_ net170 mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5847_ mod.registers.r11\[15\] _2619_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3477__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5778_ mod.registers.r10\[4\] _2580_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5734__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3745__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4729_ _1429_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5670__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__A2 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5973__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4704__C _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6150__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4011__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4946__I _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _0254_ net42 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _2439_ _2521_ _2525_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6681_ _0185_ net114 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3893_ mod.registers.r8\[9\] _3273_ _0532_ mod.registers.r10\[9\] _0863_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5632_ _2403_ _2480_ _2482_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6602__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5563_ mod.registers.r5\[13\] _2433_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6401__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4514_ _0937_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5494_ mod.registers.r4\[14\] _2380_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4445_ _1413_ _1414_ _1313_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4376_ _1343_ _1345_ _1336_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6115_ _2782_ _2791_ _2807_ _2815_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__I mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3327_ _3171_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2743_ _2757_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5652__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6681__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__A1 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6948_ _0046_ net147 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6879_ _0380_ net151 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3935__I _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__A3 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5891__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6199__A2 _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5597__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3957__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__B1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4230_ _1152_ _1196_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4685__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _1129_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4092_ _3245_ _0714_ _1059_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5634__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_370 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ _0306_ net43 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4994_ _1899_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6733_ _0237_ net62 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ _3228_ _3233_ _0728_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4070__B1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6664_ _0168_ net128 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3876_ _0631_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5615_ _2442_ _2465_ _2470_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6362__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3755__I _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _3145_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ _2422_ _2418_ _2423_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _2236_ _2367_ _2372_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4125__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4428_ _1396_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4359_ _0920_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5625__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4428__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _2743_ _2745_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__B1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6306__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout41 net44 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net54 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4600__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout63 net64 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout85 net87 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout96 net99 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_127_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4364__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__B2 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4667__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3614__B _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3875__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5616__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3627__B1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5092__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _3185_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3575__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3661_ _0415_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5400_ mod.registers.r2\[12\] _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6380_ _2952_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3592_ _3268_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _2163_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__A1 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _2172_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5855__A1 mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _0099_ net205 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4213_ _1128_ _1151_ _1167_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ _2142_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3866__B1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ _3215_ _1113_ mod.registers.r11\[9\] _1013_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3618__B1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4075_ mod.funct3\[1\] _1024_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout50_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _1944_ _1897_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6716_ _0220_ net113 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4594__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3928_ _0720_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6647_ _0151_ net127 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ mod.registers.r8\[10\] _0729_ _0730_ mod.registers.r10\[10\] _0829_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6335__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6578_ mod.des.des_counter\[2\] _2071_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_152_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4897__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _2228_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5846__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4649__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout220 net221 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4265__B _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4821__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3388__A2 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__I _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5837__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__I mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4954__I _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout185_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6262__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ mod.ldr_hzd\[11\] _1852_ _1854_ mod.ldr_hzd\[9\] _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5880_ _2556_ _2640_ _2644_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4831_ net14 _1798_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6390__B _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3379__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4576__B2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1227_ _1485_ _1369_ _1229_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6501_ mod.des.des_dout\[11\] net9 _3085_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _0556_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4693_ _1660_ _1661_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_146_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _1852_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ _0456_ _3235_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _0669_ _2714_ _2998_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3575_ _0430_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5314_ _2238_ _2254_ _2255_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6294_ _2952_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5176_ mod.pc0\[13\] _1892_ _1901_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__I _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ _1032_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__C _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4058_ _0540_ _0543_ _0546_ _0549_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5695__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3790__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6615__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4098__A3 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6765__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6906__D _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4723__B _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6547__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout100_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _3172_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5030_ mod.pc_2\[5\] _1991_ _1994_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _0079_ net105 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4246__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ mod.registers.r13\[14\] _2674_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4797__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4797__B2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5863_ _2626_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4633__B _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _1390_ _1393_ _1777_ _1780_ _1783_ _1391_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XANTENNA__4549__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5794_ mod.registers.r10\[11\] _2586_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5210__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4745_ _1030_ _1670_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6638__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3772__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4676_ _1604_ _1621_ _1627_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6415_ mod.rd_3\[3\] _2858_ _2140_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3627_ mod.registers.r3\[2\] _3165_ _0596_ mod.registers.r7\[2\] _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3763__I _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput29 net29 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3524__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6346_ _0616_ _2982_ _2986_ mod.instr\[16\] _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3558_ _0464_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6788__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ net13 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3489_ _0457_ _3259_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5277__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ mod.pc0\[12\] _1891_ _1900_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4788__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A2 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4712__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__C _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4228__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__C2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout148_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ _1474_ _1475_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _1238_ _1429_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_144_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3583__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6200_ _2102_ _2876_ _2882_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3412_ _3264_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4392_ _0789_ _0813_ _0814_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6131_ _2826_ _2827_ _2829_ _2817_ _2773_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _3193_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6062_ _2768_ _2769_ mod.pc\[0\] _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _1934_ _1912_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5303__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6964_ _0062_ net212 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5431__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _2413_ _2661_ _2666_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6895_ _0396_ net170 mod.instr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3758__I _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ _2566_ _2618_ _2622_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5195__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _2573_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3745__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _1435_ _1489_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4810__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _1353_ _1525_ _0496_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6329_ _1805_ _2975_ _2972_ mod.instr\[10\] _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_1_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5670__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__B1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6953__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5883__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5110__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3672__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3228_ _3240_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3578__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ mod.registers.r8\[14\] _2522_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ _0184_ net95 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3892_ mod.pc_2\[9\] _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5177__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5631_ mod.registers.r7\[4\] _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4924__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4630__C _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4513_ _1473_ _1482_ _1340_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ _2284_ _2379_ _2382_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4444_ _1357_ _0840_ _0875_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _1344_ _0527_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6429__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _2016_ _2809_ _2032_ _2813_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ mod.registers.r4\[0\] _3174_ _3178_ mod.registers.r1\[0\] _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _2746_ mod.pc0\[10\] _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6826__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A3 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__C _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3488__I _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4093__B _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6947_ _0045_ net147 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6878_ _0379_ net153 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5168__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5829_ _2598_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4391__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5643__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3654__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3957__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6849__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4160_ mod.registers.r14\[8\] _0891_ _0889_ mod.registers.r13\[8\] _1130_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3893__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3893__B2 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _0804_ _0806_ _0650_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_360 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_371 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _0305_ net73 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4993_ _1890_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4445__I0 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _0236_ net113 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3944_ mod.funct3\[0\] _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4070__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4070__B2 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6663_ _0167_ net132 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3875_ mod.registers.r7\[8\] _0442_ _3287_ mod.registers.r6\[8\] _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5614_ mod.registers.r6\[15\] _2466_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6412__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ net4 mod.des.des_dout\[32\] _3142_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5545_ mod.registers.r5\[9\] _2419_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3581__B1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ mod.registers.r4\[7\] _2368_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4125__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4427_ _0945_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3771__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6287__C _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A3 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4358_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3884__B2 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ mod.instr_2\[16\] _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _1248_ _1255_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5625__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _2734_ mod.pc0\[5\] _2744_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7004__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3636__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3636__B2 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3939__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4061__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout42 net44 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4600__A3 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4551__B _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout75 net83 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout86 net87 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net99 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_155_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5313__A1 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__I mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3875__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3875__B2 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5616__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3627__A1 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3627__B2 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3856__I _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout130_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3660_ mod.registers.r14\[2\] _0534_ _0535_ mod.registers.r6\[2\] _0630_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3591_ _3235_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6671__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3563__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5330_ _2238_ _2268_ _2269_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6388__B _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _2201_ _2205_ _2207_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5304__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7000_ _0098_ net209 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4212_ _1180_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5192_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3866__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3866__B2 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ _3168_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4074_ _1024_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3618__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3618__B2 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6280__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4291__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout43_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ mod.pc\[2\] _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6715_ _0219_ net111 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3766__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ mod.funct7\[1\] mod.funct7\[0\] _0617_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3397__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _0150_ net131 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3858_ _0728_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6577_ _3134_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5981__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3789_ _0458_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3554__B1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5528_ _2408_ _2404_ _2409_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3715__B _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout221 net222 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5782__A1 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3848__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3863__A4 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6227__I mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout178_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ net15 _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__B2 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5773__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _1473_ _1730_ _1340_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3586__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6500_ _3088_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3712_ _0579_ _0680_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _1495_ _1338_ _1565_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_146_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3643_ _0601_ _0604_ _0606_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6431_ _1815_ _3033_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4328__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6362_ mod.pc_1\[1\] _2995_ _2996_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3574_ _0427_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5313_ mod.registers.r1\[9\] _2246_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6293_ _2712_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ mod.des.des_dout\[23\] _2188_ _2190_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5175_ _2131_ _1925_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _1075_ _1094_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _0533_ _0536_ _0537_ _0538_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4264__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4813__C _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _1914_ _1920_ _1927_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _0133_ net126 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5216__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4120__I mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6244__A2 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4255__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4494__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _0078_ net106 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4246__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4246__B2 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _2435_ _2673_ _2676_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5994__A1 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5796__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _2538_ _2627_ _2633_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4813_ _1390_ _1776_ _1782_ _0943_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_61_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _2556_ _2585_ _2589_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4744_ _1326_ _1367_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4675_ _1572_ _1623_ _1640_ _1331_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_147_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3626_ _3169_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6414_ _3029_ _2956_ _3030_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6171__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3557_ _0460_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3524__A3 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6345_ _2985_ _2987_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6276_ mod.des.des_dout\[16\] _2933_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _3237_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _2162_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4485__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _2115_ _1925_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4109_ mod.registers.r2\[5\] _3190_ _3169_ mod.registers.r7\[5\] _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5089_ _2050_ _1896_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5985__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6732__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6882__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5976__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__B _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__B1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4460_ _1237_ _1225_ _1230_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6153__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3411_ _3236_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5900__A1 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _1352_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4703__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6130_ _2828_ _2827_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3342_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3911__B1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6396__B _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1788_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _1970_ _1976_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5967__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6963_ _0061_ net208 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ mod.registers.r13\[7\] _2662_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6605__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3978__B1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6894_ _0395_ net172 mod.instr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5719__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ mod.registers.r11\[14\] _2619_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ _2571_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4727_ _1647_ _1674_ _1685_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6144__A1 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _1320_ _1354_ _1406_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3609_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4589_ _1528_ _1529_ _1342_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _2971_ _2976_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4170__A3 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6259_ mod.instr\[12\] _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__C _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5958__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6060__I _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6438__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6628__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout160_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ _3248_ _0914_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4621__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3891_ _0552_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _2474_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6374__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4924__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5561_ _2283_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3594__I mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6126__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4512_ _1307_ _1480_ _1481_ _1337_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5492_ mod.registers.r4\[13\] _2380_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4137__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _0554_ _0860_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4688__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4374_ _0625_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6113_ _2808_ _2810_ _2032_ _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3325_ _3177_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6429__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _2722_ _2084_ _2087_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout73_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _0044_ net78 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5984__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ _0378_ net156 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5828_ _2548_ _2606_ _2611_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6365__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5168__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5759_ _2566_ _2561_ _2567_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4679__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6920__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__C1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__A2 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6356__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__B2 mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6108__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4390__I0 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _0723_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_350 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_361 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_372 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6800_ _0304_ net65 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4992_ _1934_ _1788_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_63_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6731_ _0235_ net112 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3943_ _0726_ _0810_ _0877_ _0901_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_16_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4070__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6662_ _0166_ net128 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3874_ mod.registers.r4\[8\] _0420_ _0435_ mod.registers.r15\[8\] _0844_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _2439_ _2465_ _2469_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _3144_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3581__B2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5475_ _2229_ _2367_ _2371_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4426_ _1237_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5322__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4676__A4 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5044__I mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4357_ _0716_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3308_ mod.instr_2\[17\] _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4288_ _1033_ _1256_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5979__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5086__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6943__CLK net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6027_ _2736_ _1998_ _2001_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _0027_ net202 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4061__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout43 net44 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net56 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6338__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6338__B2 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout76 net79 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_155_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5010__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6510__A1 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3324__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3627__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4824__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4052__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__B2 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ _3234_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3563__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3563__B2 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__B1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ mod.registers.r1\[4\] _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6966__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _0825_ _1177_ _1179_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5191_ mod.ins_ldr_3 mod.valid_out3 net15 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_96_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3866__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ mod.registers.r2\[9\] _0701_ _3178_ mod.registers.r1\[9\] _0596_ mod.registers.r7\[9\]
+ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _0489_ _1037_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_55_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3618__A2 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4291__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _1934_ _1912_ _1942_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6714_ _0218_ net96 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3926_ _3253_ _0886_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6645_ _0149_ net130 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3857_ _0813_ _0814_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ mod.des.des_dout\[25\] net10 _3118_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3788_ mod.pc_2\[13\] _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_118_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3554__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__I mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ mod.registers.r5\[5\] _2405_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3554__B2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3782__I _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _2358_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout200 net201 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4409_ _0950_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _2303_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout211 net212 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout222 net1 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5059__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4282__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__A2 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6839__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5782__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3793__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__CLK net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3848__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4737__B _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__I _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5470__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4025__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4760_ _1665_ _1535_ _1729_ _1422_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3711_ _3261_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4691_ _1420_ _1568_ _1569_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6430_ _3040_ _3042_ _3023_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3642_ mod.registers.r14\[2\] _0607_ _0608_ mod.registers.r13\[2\] _0611_ _0612_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _3263_ _2714_ _2997_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3573_ mod.registers.r13\[7\] _0541_ _0542_ mod.registers.r1\[7\] _0543_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6292_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__A1 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5243_ _0628_ _2191_ _2174_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ mod.pc\[13\] _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ _0899_ _0574_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_96_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ _0458_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5461__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4264__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3777__I mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _1921_ _1922_ _1923_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3909_ _3170_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5992__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ mod.ldr_hzd\[0\] _1856_ _1858_ mod.ldr_hzd\[2\] mod.instr_2\[5\] _1859_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6628_ _0132_ net76 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4319__A3 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ mod.des.des_dout\[17\] net2 _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout190_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ mod.registers.r13\[13\] _2674_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5994__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5861_ mod.registers.r12\[3\] _2629_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4812_ _1781_ _1394_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5792_ mod.registers.r10\[10\] _2586_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4743_ _1708_ _1711_ _1712_ _1332_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4674_ _1366_ _1641_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3509__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6413_ mod.rd_3\[2\] _2858_ _2140_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3625_ _0489_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6171__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _0480_ _2982_ _2986_ mod.instr\[15\] _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3556_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6275_ mod.instr\[16\] _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3487_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5157_ mod.pc\[12\] _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6684__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3693__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ _1024_ _3259_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5088_ mod.pc\[8\] _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5987__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4891__I mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4039_ mod.registers.r12\[7\] _0888_ _0608_ mod.registers.r13\[7\] _1009_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5227__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3515__A4 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3920__B2 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5673__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__I _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3684__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5976__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3739__B2 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout203_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3410_ mod.pc_2\[0\] _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__4164__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1355_ _1359_ _0497_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4976__I mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3911__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3341_ _3193_ _3162_ _3182_ _3184_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1389_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ _1794_ _1968_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5416__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4219__A2 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3427__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6962_ _0060_ net208 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5967__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _2410_ _2661_ _2665_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3978__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6893_ _0394_ net172 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _2564_ _2618_ _2621_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5775_ _2538_ _2572_ _2578_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4726_ _3242_ _1680_ _1691_ _1659_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_147_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4657_ _1301_ _1623_ _1626_ _1432_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4155__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3608_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4588_ _1556_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_150_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3902__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _1781_ _2975_ _2972_ mod.instr\[9\] _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3539_ mod.registers.r4\[6\] _0508_ _3237_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _2924_ _2925_ _2926_ _2917_ _2923_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4458__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6189_ _2033_ _2868_ _2875_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3965__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4394__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3406__S _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5646__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout153_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3890_ _0813_ _0814_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6251__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _2431_ _2432_ _2434_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4511_ _1351_ _1336_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6126__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5491_ _2276_ _2379_ _2381_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4137__A1 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4137__B2 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _0627_ _1410_ _1411_ _1333_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5885__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4373_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4639__C _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6112_ _2802_ _1885_ mod.pc\[7\] _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3324_ _3175_ _3176_ _3163_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6429__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5637__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6043_ _2730_ _2069_ _2755_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6722__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6945_ _0043_ net77 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _0377_ net155 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__B1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5827_ mod.registers.r11\[7\] _2607_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6365__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ mod.registers.r9\[14\] _2562_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4709_ _1442_ _1254_ _1513_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5689_ _2422_ _2515_ _2518_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4128__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__B _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6053__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__B1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__A1 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__C2 _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3811__B1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6356__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6600__I0 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5867__A1 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_340 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_351 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_362 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_373 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _1915_ _1950_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6730_ _0234_ net97 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6895__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3942_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3802__B1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _0165_ net129 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3873_ mod.pc_2\[8\] _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5612_ mod.registers.r6\[14\] _2466_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6592_ net3 mod.des.des_dout\[31\] _3142_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5543_ _2253_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5474_ mod.registers.r4\[6\] _2368_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4425_ _0992_ _1394_ _1391_ _1379_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3869__B1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _1307_ _1314_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3307_ _3158_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _0551_ _1022_ _1026_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5086__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4833__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6156__I _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4597__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _0026_ net186 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout44 net46 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6859_ _0360_ net191 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout66 net67 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout77 net78 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout88 net89 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout99 net100 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5010__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6618__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6768__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A2 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6274__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4588__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A3 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6015__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5001__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout116_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3563__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4760__B2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4210_ _1177_ _1179_ _0826_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4512__B2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1861_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4141_ mod.registers.r12\[9\] _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _1038_ _1039_ _1040_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_96_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ _1915_ _1933_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6713_ _0217_ net111 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3925_ _0890_ _0892_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _0148_ net79 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _3133_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4200__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3787_ _0728_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5526_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3554__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5457_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4408_ _0987_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout201 net202 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5388_ _2301_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout212 net222 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3857__A3 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _0454_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5059__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6009_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3490__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A3 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4134__I _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3793__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5470__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _0669_ _0528_ _0674_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4981__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _1339_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3641_ _0609_ _3213_ _3214_ _3218_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6933__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ mod.pc_1\[0\] _2995_ _2996_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3572_ _0448_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ mod.des.des_dout\[30\] _2248_ _2250_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ mod.valid1 _2709_ _2151_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_114_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5289__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ _2169_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _2092_ _2122_ _2129_ _1896_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ _1076_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6238__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4055_ _3226_ _0618_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4663__B _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__A1 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4957_ mod.pc\[1\] _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3908_ _0799_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4972__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _0131_ net74 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3839_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4724__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _3118_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ mod.registers.r5\[1\] _2391_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6489_ _3082_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4129__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6806__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3968__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4963__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4191__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5691__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout183_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5994__A3 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5860_ _2536_ _2627_ _2632_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4811_ _0942_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _2554_ _2585_ _2588_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _1346_ _1335_ _1400_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4673_ _1072_ _1549_ _1642_ _1060_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6203__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _2141_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3624_ _0576_ _0592_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4706__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6343_ _2950_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3555_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6459__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6459__B2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6274_ _2936_ _2937_ _2938_ _2929_ _2935_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3486_ _3234_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4658__B _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5225_ mod.des.des_dout\[21\] _2167_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5131__A1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6829__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _2092_ _2108_ _2113_ _1924_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_29_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3693__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__B2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ mod.funct3\[0\] _1023_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _2041_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4038_ _1005_ _1006_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6979__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5198__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _2712_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6113__B _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__I _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__A1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5122__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5673__A2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3684__B2 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__I _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4936__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4750__C _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__C1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5361__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3340_ mod.instr_2\[17\] _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3911__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _1971_ _1972_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3675__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5416__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3427__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6961_ _0059_ net208 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3427__B2 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__B _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5912_ mod.registers.r13\[6\] _2662_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3401__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3978__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _0393_ net172 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5843_ mod.registers.r11\[13\] _2619_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ mod.registers.r10\[3\] _2574_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4725_ _0922_ _1408_ _1693_ _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5328__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4232__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4656_ _1495_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3607_ _3265_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5352__A1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _1401_ _0912_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6651__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3538_ _0418_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6326_ _2955_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5104__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ mod.des.des_dout\[11\] _2921_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3469_ _3284_ _0416_ _0425_ _0426_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _1850_ _2143_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7007__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6188_ mod.pc_1\[7\] _2869_ _2873_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _2095_ _2097_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5407__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6080__A2 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4407__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3969__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4091__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5591__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4394__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4146__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A1 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3981__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5646__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__A4 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout146_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5582__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6674__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4510_ _0776_ _0803_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ mod.registers.r4\[12\] _2380_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4137__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _0790_ _0775_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3891__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4372_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3896__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _2017_ _2780_ _2812_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3323_ mod.instr_2\[14\] _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6042_ _2729_ mod.pc0\[9\] _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5637__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__I0 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3840__B _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout59_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6062__A2 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _0042_ net152 mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4073__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6875_ _0376_ net180 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3820__B2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5826_ _2546_ _2606_ _2610_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5573__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _2289_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _1675_ _1676_ _1440_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5688_ mod.registers.r8\[9\] _2516_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5325__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4128__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _1468_ _0555_ _1608_ _0623_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ mod.instr_2\[3\] _2958_ _2963_ mod.instr\[3\] _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3306__I mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4300__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4064__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4064__B2 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__B2 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6697__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6600__I1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4756__B _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_330 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_341 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_352 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_363 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_374 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _1952_ _1955_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _0908_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3802__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3802__B2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3872_ _0812_ _0827_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6660_ _0164_ net77 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ _2436_ _2465_ _2468_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6591_ _3143_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3566__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5542_ _2417_ _2418_ _2420_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4763__C1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5307__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _2218_ _2367_ _2370_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5606__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__B1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4424_ _1376_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__B2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ _1315_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3306_ mod.instr_2\[14\] _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ mod.pc_2\[6\] _1205_ _0510_ _0523_ _1047_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_86_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4294__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4046__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6927_ _0025_ net186 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5794__A1 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3796__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6858_ _0359_ net190 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout45 net46 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout56 net66 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout67 net89 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5809_ _2597_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5546__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4349__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout78 net79 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout89 net146 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6594__I0 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _0293_ net103 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__I _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4420__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A3 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5251__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4037__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__B2 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6082__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__I0 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4330__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4140_ _0888_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6265__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ mod.registers.r12\[6\] _0887_ _3211_ mod.registers.r13\[6\] _1041_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6862__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4028__B2 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _1916_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6712_ _0216_ net95 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3924_ mod.registers.r2\[4\] _0893_ _3174_ mod.registers.r4\[4\] mod.registers.r10\[4\]
+ _0602_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5528__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ _0147_ net76 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6576__I0 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3855_ mod.pc_2\[11\] _0777_ _0819_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6574_ mod.des.des_dout\[24\] net9 _3129_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4200__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3786_ _0683_ _0684_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4200__B2 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _2217_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5456_ _2358_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5700__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5387_ _2236_ _2309_ _2314_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout202 net203 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_132_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout213 net215 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4338_ _0683_ _0684_ _0680_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4269_ _0988_ _0990_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6008_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A3 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3490__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5020__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__I _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6885__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3481__A2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ mod.registers.r15\[2\] _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6183__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _0446_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4733__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5310_ _2213_ _2251_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6290_ _2948_ _2889_ _2949_ _2891_ _2742_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__I mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5241_ _2136_ _1604_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _2126_ _2127_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4123_ _3238_ _1078_ _1088_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6238__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4054_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput2 io_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6608__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout41_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4956_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6758__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3907_ _0811_ _0842_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4972__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4887_ _1849_ mod.instr_2\[3\] _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6174__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _0130_ net71 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3838_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4185__B1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _3123_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5921__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ mod.registers.r4\[12\] _0738_ _3266_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6488_ mod.des.des_dout\[5\] net3 _3080_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _2261_ _2343_ _2347_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4488__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3314__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__C2 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6561__S _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4191__A3 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5704__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout176_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4483__C _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6900__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ _1390_ _1778_ _1779_ _1392_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ mod.registers.r10\[9\] _2586_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4403__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _1328_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _1072_ _0944_ _0938_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _1849_ _2883_ _3028_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5903__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3509__A3 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3623_ _0495_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6342_ _2707_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3554_ mod.pc_2\[6\] _0499_ _0510_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6273_ mod.des.des_dout\[15\] _2933_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3485_ _3254_ _3180_ _3222_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_103_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _3263_ _2168_ _2170_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5131__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout89_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _2092_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3693__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4106_ _0591_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_96_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5086_ _1970_ _2040_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_57_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ mod.registers.r11\[7\] _0605_ _3199_ mod.registers.r9\[7\] _1007_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _2711_ _1884_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4939_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _0113_ net85 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3309__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5370__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6556__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4881__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6923__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4633__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4149__B1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__C2 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A3 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6310__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3675__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3889__I _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6960_ _0058_ net213 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3427__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ _2407_ _2661_ _2664_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6891_ _0392_ net172 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ _2560_ _2618_ _2620_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5773_ _2536_ _2572_ _2577_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4724_ _0526_ _1103_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4655_ _1260_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3606_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4586_ _1555_ _0454_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6325_ _2971_ _2974_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3537_ mod.registers.r11\[6\] _0505_ _0506_ mod.registers.r2\[6\] _0507_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_143_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _2718_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5104__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3468_ mod.registers.r15\[0\] _0435_ _0437_ mod.registers.r12\[0\] _0438_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ mod.rd_3\[0\] _2144_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _2017_ _2868_ _2874_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A1 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3399_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5138_ _0957_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5069_ _1911_ _2004_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4615__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3969__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__A1 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3748__B _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5591__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4394__A3 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A3 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3354__A1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5254__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4298__C _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4606__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4082__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4909__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6819__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout139_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4440_ _1409_ _0827_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6531__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3345__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4371_ _0621_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3896__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6110_ _2767_ _2811_ _2778_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ mod.instr_2\[15\] _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__I1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3412__I _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _0041_ net154 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4073__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6874_ _0375_ net178 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3820__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3568__B _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ mod.registers.r11\[6\] _2607_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _2564_ _2561_ _2565_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5573__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3584__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _1515_ _1252_ _1249_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5687_ _2417_ _2515_ _2517_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6522__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _1316_ _0576_ _0592_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4569_ _1538_ _0724_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6308_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5089__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ mod.instr\[7\] _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4836__A1 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3322__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5564__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__I _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5316__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3327__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3878__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_320 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_331 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_342 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_353 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_364 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_375 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3940_ _3227_ _0902_ _0909_ _0903_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3802__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3871_ _0828_ _0553_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5610_ mod.registers.r6\[13\] _2466_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6590_ net2 mod.des.des_dout\[30\] _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3566__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3566__B2 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5541_ mod.registers.r5\[8\] _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4763__B1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4763__C2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ mod.registers.r4\[5\] _2368_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5307__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3318__A1 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__B2 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4423_ _1391_ _1380_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _1317_ _1319_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ mod.instr_2\[15\] _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4285_ _1249_ _1252_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6024_ _2706_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout71_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A1 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4046__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _0024_ net187 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _0358_ net191 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout46 net67 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout57 net61 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout68 net72 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout79 net82 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5546__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _0292_ net68 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4349__A3 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6594__I1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5739_ _2550_ _2551_ _2553_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3317__I _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5482__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4285__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__I1 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5707__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3720__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6538__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4070_ mod.registers.r14\[6\] _3208_ _3169_ mod.registers.r7\[6\] _1040_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5473__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4028__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__A1 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4972_ _1051_ _1935_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _0215_ net96 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5110__C _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3923_ _3191_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6642_ _0146_ net70 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5528__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3854_ _0820_ _0821_ _0822_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6576__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3539__A1 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _3132_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5617__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3785_ _0727_ _0728_ _0740_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4200__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ _2403_ _2404_ _2406_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _2356_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4406_ _1245_ _1247_ _1303_ _1304_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_132_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5161__B1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5700__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ mod.registers.r2\[7\] _2310_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout203 net204 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4337_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6687__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4268_ _1225_ _1230_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5464__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _2711_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4806__A4 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ mod.registers.r11\[11\] _0705_ _0697_ mod.registers.r1\[11\] _1169_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _0007_ net149 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6192__A2 _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6559__S _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6358__I _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3702__B2 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5455__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5207__A1 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3510__I _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout121_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout219_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3570_ mod.registers.r15\[7\] _0435_ _0437_ mod.registers.r12\[7\] _0540_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5930__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _2182_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _2126_ _2127_ _2056_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _0615_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4249__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4053_ _3232_ _3251_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_84_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__I _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _1895_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _0802_ _0860_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4886_ mod.instr_2\[4\] mod.instr_2\[3\] _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _0129_ net85 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3837_ _0804_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6174__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4185__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ mod.des.des_dout\[16\] net19 _3119_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4185__B2 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5921__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3768_ _0419_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5507_ _2185_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6487_ _3081_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3699_ mod.pc_2\[1\] _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_105_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ mod.registers.r3\[10\] _2344_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4488__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5369_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5810__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__B2 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6702__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6852__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5912__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3518__A4 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5428__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4100__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4336__I _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout169_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _1352_ _1630_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3611__B1 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ _1315_ _1314_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4167__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ mod.rd_3\[1\] _2884_ _3017_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3622_ _0579_ _0591_ _3262_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6341_ _2978_ _2984_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3553_ _0513_ _0516_ _0519_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_155_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _2718_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3484_ _3246_ _3262_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5667__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3678__B1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ mod.pc_2\[12\] _1089_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_96_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5419__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3693__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4105_ _0578_ _1074_ _0896_ _0898_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__5630__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ _1970_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6092__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4036_ mod.registers.r2\[7\] _0701_ _3195_ mod.registers.r10\[7\] _1006_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ net12 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6395__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4938_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4869_ _1814_ _1835_ _1015_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _0112_ net86 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3905__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _3094_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5658__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5540__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4584__C _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4633__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6138__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__B2 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5715__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__C1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4321__B2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A1 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ mod.registers.r13\[5\] _2662_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6898__CLK net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6890_ _0391_ net170 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5841_ mod.registers.r11\[12\] _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4388__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ mod.registers.r10\[2\] _2574_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4723_ _1675_ _1669_ _1484_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_147_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _1071_ _1267_ _1056_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5888__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3605_ _0556_ _0557_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4585_ _1265_ _1070_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3899__B1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _1391_ _2968_ _2972_ mod.instr\[8\] _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3536_ _0411_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4560__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ mod.instr\[11\] _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3467_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5206_ _1849_ _2143_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4312__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6186_ mod.pc_1\[6\] _2869_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3398_ _3230_ _3231_ mod.instr_2\[1\] _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4863__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5137_ mod.funct7\[0\] _1206_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6065__A1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _2005_ _2024_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5812__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4615__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4019_ _0799_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5879__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3339__C1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4146__A4 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3354__A2 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4303__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6366__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A3 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3593__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6531__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout201_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ _3173_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6040_ _2752_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__C1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5180__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6942_ _0040_ net152 mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__A3 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6873_ _0374_ net177 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5824_ _2544_ _2606_ _2609_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ mod.registers.r9\[13\] _2562_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3584__A2 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _0526_ _1103_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5686_ mod.registers.r8\[8\] _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ _1572_ _1605_ _1606_ _1515_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4568_ _0899_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3519_ _3252_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6307_ _2950_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4499_ _1468_ _1305_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6286__A1 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6238_ _2908_ _2901_ _2910_ _2905_ _2911_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4836__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _1893_ _2859_ _2862_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6038__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4049__B1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5261__A2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3732__C1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_310 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6029__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_321 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_332 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_343 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_354 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_365 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_376 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6936__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ _2390_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3566__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _2205_ _2367_ _2369_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3318__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _0914_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4353_ _1317_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3304_ _3157_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ _1253_ _1093_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _2739_ _2740_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3423__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4046__A3 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ _0023_ net195 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6856_ _0357_ net192 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout47 net51 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout58 net61 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5807_ _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4203__B1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout69 net72 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3999_ mod.registers.r6\[15\] _0966_ _0967_ mod.registers.r5\[15\] _0968_ mod.registers.r8\[15\]
+ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6787_ _0291_ net68 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ mod.registers.r9\[8\] _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5669_ _2394_ _2502_ _2506_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3333__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3493__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6431__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3489__B _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3508__I _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3484__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _1917_ _1937_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6710_ _0214_ net90 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6490__S _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3922_ mod.registers.r14\[4\] _0891_ _0705_ mod.registers.r11\[4\] _0892_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3853_ mod.registers.r13\[11\] _0520_ _0521_ mod.registers.r1\[11\] _0823_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6641_ _0145_ net85 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3539__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3784_ _0742_ _0744_ _0750_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6572_ mod.des.des_dout\[23\] net8 _3129_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ mod.registers.r5\[4\] _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5454_ _2155_ _2157_ _2159_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3862__B _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4405_ _1326_ _1330_ _1348_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5161__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5385_ _2229_ _2309_ _2313_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5161__B2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout204 mod.clk net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4336_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout215 net216 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4267_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6006_ _2724_ _2727_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5464__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4198_ mod.registers.r14\[11\] _0891_ _0703_ mod.registers.r9\[11\] mod.registers.r2\[11\]
+ _0893_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6413__A1 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6908_ _0409_ net161 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _0340_ net177 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5808__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__B _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3328__I _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3702__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6781__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3466__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3998__I _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3769__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5718__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4718__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__I _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ mod.pc_2\[13\] _0955_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _1089_ _1090_ _0617_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4052_ _3254_ _1008_ _1020_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_37_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3457__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 io_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_110_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4957__A1 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _1900_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3905_ _0828_ _0861_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4885_ mod.ldr_hzd\[3\] _1852_ _1854_ mod.ldr_hzd\[1\] _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6624_ _0128_ net87 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3836_ _0577_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4185__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5382__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _3122_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3767_ mod.registers.r11\[12\] _0735_ _0736_ mod.registers.r2\[12\] _0737_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6654__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5506_ _2386_ _2389_ _2392_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3698_ _0650_ _0666_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6486_ mod.des.des_dout\[4\] net2 _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5437_ _2254_ _2343_ _2346_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ _2300_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3696__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3696__B2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _0731_ _0734_ _0737_ _0739_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5299_ _1951_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5538__I _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5373__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4598__B _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3687__A1 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4100__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3611__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _1420_ _1632_ _1634_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _0580_ _0421_ _0585_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5364__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ mod.registers.r13\[6\] _0520_ _0521_ mod.registers.r1\[6\] _0522_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6340_ _1136_ _2982_ _2979_ mod.instr\[14\] _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6271_ mod.instr\[15\] _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6279__I mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5116__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3483_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4301__B _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5667__A2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5222_ _2171_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3678__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3678__B2 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4875__C2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _2094_ _2098_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5419__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4104_ _0567_ _0572_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _0843_ _2042_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6092__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4035_ mod.registers.r15\[7\] _0963_ _3186_ mod.registers.r6\[7\] _3189_ mod.registers.r5\[7\]
+ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3850__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__B2 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ mod.valid0 _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ mod.des.des_counter\[0\] _3150_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _1833_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5355__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _0111_ net159 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3819_ _0784_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _1665_ _1360_ _1367_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6538_ _3092_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3905__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__B1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3606__I _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _1819_ _3064_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3669__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__A1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__I _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__B1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__C2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4321__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout181_I net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4347__I _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4085__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4624__A3 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _2600_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4388__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _2534_ _2572_ _2576_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3596__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4722_ _1675_ _1670_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4653_ _1445_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5906__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3604_ _0567_ _0572_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4584_ _1517_ _1522_ _1523_ _1553_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__B2 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__C _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6323_ _2971_ _2973_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3535_ _3290_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3426__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _2920_ _2913_ _2922_ _2917_ _2923_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_fanout94_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3466_ _3281_ _0417_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5205_ mod.rd_3\[1\] _2144_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4312__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3397_ _3244_ _3247_ _3249_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_69_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5136_ mod.pc_2\[11\] _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5067_ _1790_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6842__CLK net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4018_ _0950_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3823__B2 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A2 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2680_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3339__B1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3339__C2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__I0 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3336__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4303__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A2 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A4 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5319__A1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3593__A3 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5726__I _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6715__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3345__A3 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3320_ _3166_ _3168_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6295__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6865__CLK net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3502__B1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__C2 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4058__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _0039_ net154 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3805__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6872_ _0373_ net187 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5823_ mod.registers.r11\[5\] _2607_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ _2283_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4705_ _0526_ _1103_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3584__A3 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ _2503_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _1454_ _1448_ _1453_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5730__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _1401_ _0623_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6306_ _2759_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3518_ _0472_ _0474_ _0475_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _0691_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _2788_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3449_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ mod.pc_1\[0\] _2861_ _2822_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__A2 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _2060_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4049__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6099_ _1389_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4049__B2 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5013__A3 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3732__B1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__C2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_300 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_311 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_322 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_333 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_344 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_355 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_366 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_377 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5788__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3799__B1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout144_I net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5456__I _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__B1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5470_ mod.registers.r4\[4\] _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ _3229_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6488__S _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4352_ _1320_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_140_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6268__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3303_ mod.des.des_counter\[2\] _3151_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4283_ _0591_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6022_ _2726_ _1983_ _2731_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout57_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6924_ _0022_ net197 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6855_ _0356_ net192 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5806_ _2327_ _2499_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout48 net51 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout59 net61 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4203__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _0290_ net68 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4203__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3998_ _0473_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5737_ _2531_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5951__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__I _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ mod.registers.r8\[1\] _2504_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5703__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _0938_ _1588_ _1061_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5599_ _2417_ _2459_ _2461_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__B2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5942__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4745__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3705__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5170__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5225__B _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__CLK net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ _1206_ _0492_ _1045_ _0669_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__4433__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _3208_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6640_ _0144_ net129 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3852_ mod.registers.r5\[11\] _0517_ _0518_ mod.registers.r7\[11\] _0822_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4736__A2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _3131_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5186__I _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ mod.registers.r9\[12\] _0751_ _0752_ mod.registers.r3\[12\] _0753_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5522_ _2390_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5453_ _2355_ _2149_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4404_ _0992_ _1349_ _1361_ _1368_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5384_ mod.registers.r2\[6\] _2310_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5161__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _0808_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout205 net207 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3434__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout216 net221 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4266_ _1004_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _2726_ _1903_ _0003_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4197_ _1165_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6413__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _0408_ net160 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _0339_ net181 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4188__B1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5924__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4727__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _0273_ net73 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3609__I _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5152__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3344__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3466__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4663__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3519__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__B2 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ mod.funct7\[1\] _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4051_ _3264_ _1002_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_36_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__B2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4957__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4953_ _1890_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4884_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__C _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6623_ _0127_ net161 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3835_ _0560_ _0618_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6554_ mod.des.des_dout\[15\] net18 _3119_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3766_ _0412_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5382__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ mod.registers.r5\[0\] _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ _3074_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3697_ _0528_ _0552_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_106_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ mod.registers.r3\[9\] _2344_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5134__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6949__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5367_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3696__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4893__A1 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4318_ _1226_ _1202_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5298_ _2208_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ _1152_ _1218_ _1143_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4645__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5819__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5373__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6322__B2 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3687__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6086__B1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6389__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5729__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A2 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _0586_ _0587_ _0588_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4167__A3 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3551_ _0448_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6270_ _2932_ _2925_ _2934_ _2929_ _2935_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5116__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ _3263_ _3266_ _0423_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_142_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4175__I0 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5221_ _1792_ _3257_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3678__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4875__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__B2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5152_ mod.pc_2\[11\] _2097_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _1056_ _1060_ _1064_ _1071_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_57_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _2043_ _2028_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4034_ _0779_ _1003_ _0789_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _1895_ _1884_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5639__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4936_ _3224_ _1905_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _1820_ _1834_ _1835_ _1819_ _1836_ _1818_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_20_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6606_ _0110_ net84 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3818_ _0785_ _0786_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5355__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _1352_ _1324_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6537_ _2427_ _3106_ _3111_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3905__A3 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3749_ _0595_ _0699_ _0710_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5107__A2 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _3068_ _3069_ _3057_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6304__B2 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5419_ _2194_ _2330_ _2335_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ net20 _2152_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3669__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4094__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__A1 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__A1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__B _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3357__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5284__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4857__B2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3532__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout174_I net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6644__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A4 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ mod.registers.r10\[1\] _2574_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3596__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6794__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _1689_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3596__B2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6534__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ _1580_ _1261_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3348__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3603_ mod.pc_2\[4\] _0499_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4583_ _1331_ _1543_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4312__B _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6322_ _1392_ _2968_ _2972_ mod.instr\[7\] _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3534_ mod.registers.r14\[6\] _0502_ _0503_ mod.registers.r6\[6\] _0504_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4560__A3 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6253_ _2741_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3465_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6184_ _2752_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout87_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _3248_ _3228_ mod.funct3\[0\] _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_97_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _2093_ _2080_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3442__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ mod.pc_2\[7\] _2025_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5273__A1 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4017_ _3247_ _0958_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3823__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _2427_ _2694_ _2699_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _1885_ _1887_ mod.valid0 _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5899_ _2385_ _2654_ _2657_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6525__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3339__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3339__B2 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__I1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4839__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3511__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6667__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5016__B2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__C1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3527__I _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3345__A4 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4358__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3502__B2 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5255__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _0038_ net162 mod.rd_3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3805__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6871_ _0372_ net186 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5189__I _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _2540_ _2606_ _2608_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3569__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _2560_ _2561_ _2563_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5917__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4230__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _1654_ _1657_ _1658_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ _2501_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _1300_ _0940_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1501_ _1419_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5730__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _2760_ _2960_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3517_ _0479_ _0481_ _0484_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_89_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4497_ _0726_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6236_ mod.des.des_dout\[6\] _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3448_ _0415_ _0416_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4297__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6167_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _3230_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5118_ _2059_ _2061_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6098_ _2783_ _2791_ _2798_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4049__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__A1 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5049_ _2008_ _2009_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_38_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3980__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5182__B1 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3732__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3732__B2 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__I _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4288__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4532__I0 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_301 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_312 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_323 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_334 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_345 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5237__A1 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_356 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_367 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_378 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3799__A1 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5737__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout137_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3971__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__B2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _3227_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3723__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _0579_ _0525_ _0681_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_99_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ _3156_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_125_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4282_ _1250_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _2723_ mod.pc0\[4\] _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4816__I _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _0021_ net195 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6854_ _0355_ net198 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5805_ _2568_ _2591_ _2596_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout49 net51 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6785_ _0289_ net45 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4203__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _0468_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__A1 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ _2529_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _2386_ _2502_ _2505_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4618_ _1056_ _1549_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5703__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ mod.registers.r6\[8\] _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4549_ _1518_ _1514_ _1075_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6503__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ mod.des.des_dout\[2\] _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6705__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3786__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6855__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3705__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3705__B2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4130__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3484__A3 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5241__B _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3920_ mod.registers.r12\[4\] _0888_ _0889_ mod.registers.r13\[4\] _0890_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3641__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ mod.registers.r9\[11\] _0511_ _0512_ mod.registers.r3\[11\] _0821_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6072__B _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4371__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6570_ mod.des.des_dout\[22\] net7 _3129_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3782_ _0512_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4736__A3 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _2388_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6499__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _2146_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5697__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _0990_ _1369_ _1372_ _1246_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5383_ _2218_ _2309_ _2312_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4334_ _1298_ _1299_ _3241_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout206 net207 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout217 net218 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5449__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6497__I0 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4265_ _3247_ _1231_ _1232_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6004_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4196_ _1161_ _1164_ _0839_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4672__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3450__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _0407_ net161 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4975__A3 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _0338_ net177 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4281__I _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__B2 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5924__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6768_ _0272_ net57 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__A3 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5719_ mod.registers.r9\[3\] _2532_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6699_ _0203_ net111 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5688__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3625__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__I _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4360__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5840__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__I _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4179__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__A2 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3535__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ _1009_ _1018_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4406__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ mod.pc0\[1\] _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3903_ _0862_ _0464_ _0867_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6159__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ mod.instr_2\[4\] _1850_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3834_ _3253_ _0599_ _0613_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6622_ _0126_ net161 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3917__A1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _3121_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3765_ _3291_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4969__C _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6484_ _3079_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3696_ _0651_ _0464_ _0656_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5435_ _2245_ _2343_ _2345_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4893__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ _1276_ _1286_ _1223_ _1203_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ _2191_ _2040_ _2209_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _1213_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3448__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4276__I _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ _0858_ _1147_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3853__B1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6322__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5570__I _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6086__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__B1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5833__A1 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4914__I _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4167__A4 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout217_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3550_ _0446_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3481_ _0432_ _0438_ _0443_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_127_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ mod.ins_ldr_3 mod.valid_out3 net15 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4175__I1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4875__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _1987_ _2108_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4102_ _1062_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5082_ _0530_ _2025_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5824__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _0687_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2708_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _3225_ _1387_ _1903_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4866_ _1135_ _1136_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _0109_ net84 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6916__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3817_ mod.registers.r14\[14\] _0732_ _0730_ mod.registers.r10\[14\] _0787_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4012__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _1345_ _1481_ _1638_ _1467_ _1660_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4563__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6536_ mod.registers.r15\[11\] _3107_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3748_ _0624_ _0693_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3679_ _0644_ _0645_ _0646_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6467_ _3055_ _3036_ _3066_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6304__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ mod.registers.r3\[2\] _2332_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6398_ _2152_ _3020_ _2831_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3669__A3 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5349_ _2168_ _2136_ _1435_ _2273_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_87_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5815__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6435__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6170__B _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4003__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6543__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3357__A2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5806__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4609__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4085__A3 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout167_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6939__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3596__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _1467_ _1421_ _1540_ _1566_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4651_ _1607_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6534__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3602_ _0568_ _0569_ _0570_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4545__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4582_ _1367_ _1546_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3533_ _3286_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6321_ _2962_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6252_ mod.des.des_dout\[10\] _2921_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ _0429_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _3244_ _2152_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6183_ _1999_ _2868_ _2871_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3395_ _3226_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5134_ mod.pc_2\[10\] _0958_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _2026_ _2012_ _2027_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5273__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4016_ _0687_ _0984_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5025__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ mod.registers.r14\[11\] _2695_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4918_ net13 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4784__B2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5898_ mod.registers.r13\[0\] _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4849_ mod.ldr_hzd\[14\] _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3339__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _3094_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6289__A1 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__I _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3633__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3511__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3814__A3 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4224__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__C2 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5295__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3808__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3971__C _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6611__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3502__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3805__A3 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4374__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6870_ _0371_ net187 mod.pc_1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ mod.registers.r11\[4\] _2607_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3569__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4766__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ mod.registers.r9\[12\] _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4230__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ _1664_ _1668_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5683_ _2414_ _2509_ _2514_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4518__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4634_ _1585_ _1586_ _1590_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ _1532_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6304_ _0903_ _2958_ _2951_ mod.instr\[2\] _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3516_ mod.registers.r15\[1\] _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4496_ _3242_ _1461_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6235_ _2888_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3447_ _3270_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5494__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6166_ _2856_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3378_ mod.instr_2\[0\] _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _2076_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6097_ _1980_ _2766_ _2800_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6443__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ mod.pc_2\[5\] _1991_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input12_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _0097_ net209 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5182__B2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6634__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3732__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5999__B _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__C1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6784__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_302 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_313 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_324 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_335 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_346 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_357 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_368 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_379 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3799__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4922__I _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ _0757_ _0861_ _0551_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3723__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3301_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_113_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4281_ _0574_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6020_ _2708_ _2738_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6425__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _0020_ net195 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4987__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__A3 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6853_ _0354_ net199 mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ mod.registers.r10\[15\] _2592_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4739__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout39 net40 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6784_ _0288_ net43 mod.registers.r12\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _0600_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5735_ _2244_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5666_ mod.registers.r8\[0\] _2504_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4617_ _1306_ _1407_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5663__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ _2447_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _1073_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _0812_ _1069_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _2888_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3478__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__B1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6494__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _2816_ _2837_ _2841_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6416__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__B2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4130__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6407__A1 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4969__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3641__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__B2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3850_ mod.registers.r15\[11\] _0514_ _0515_ mod.registers.r12\[11\] _0820_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3781_ _0511_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5394__A1 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5520_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5146__A1 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__I _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _2296_ _2349_ _2354_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4601__B _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5697__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4402_ _0988_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ mod.registers.r2\[5\] _2310_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4333_ _1298_ _1299_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout207 net208 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout218 net220 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__6497__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4264_ _0926_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6003_ _2711_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3731__I _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ _0839_ _1161_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout62_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3880__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5621__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6905_ _0406_ net162 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6836_ _0337_ net180 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4188__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5385__A1 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _0271_ net57 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3979_ _3243_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4727__A4 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5718_ _2198_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ _0202_ net98 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5137__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5649_ _2472_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5688__A2 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__B _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3871__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4472__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5376__A1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3926__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4351__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6479__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3551__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 io_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3862__A1 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5603__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4951_ _1915_ _1910_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3614__A1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5478__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4382__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3902_ _0868_ _0869_ _0870_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4882_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4315__C _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _0125_ net159 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3833_ _0790_ _0800_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3927__S _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ mod.des.des_dout\[14\] net17 _3119_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3764_ mod.registers.r14\[12\] _0732_ _0733_ mod.registers.r6\[12\] _0734_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _2387_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6316__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6483_ mod.des.des_dout\[3\] net19 _3075_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3726__I _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _0657_ _0658_ _0659_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_106_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5434_ mod.registers.r3\[8\] _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ _2150_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4316_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5296_ mod.pc_2\[8\] _2221_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4247_ _1214_ _1215_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3461__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4178_ _0858_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3853__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3853__B2 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3605__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6995__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__B1 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _0323_ net41 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__B _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__B2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4636__A3 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5298__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__I _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6718__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout112_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3780__B1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3480_ mod.registers.r13\[0\] _0447_ _0449_ mod.registers.r1\[0\] _0450_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6868__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _2107_ _1489_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6078__B mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4101_ _1068_ _0929_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_96_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ _0530_ _2025_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__A3 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4032_ mod.funct7\[2\] _0614_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3835__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _2708_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5052__A3 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3599__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4934_ _3155_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _0480_ _3256_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6604_ _0108_ _0003_ net218 mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3816_ mod.registers.r13\[14\] _0745_ _0738_ mod.registers.r4\[14\] _0733_ mod.registers.r6\[14\]
+ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4012__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4012__B2 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1760_ _1761_ _3243_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6535_ _2424_ _3106_ _3110_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4563__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3456__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3747_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ _1818_ _3064_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3678_ mod.registers.r13\[2\] _0541_ _0542_ mod.registers.r1\[2\] _0647_ _0648_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5417_ _2186_ _2330_ _2334_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4315__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ mod.valid_out3 _2153_ _2713_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _2270_ _2284_ _2285_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3405__B _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5279_ _0902_ _0561_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4251__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4003__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4003__B2 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4554__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3366__I mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4306__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3817__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__B2 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__I _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _0918_ _1614_ _1615_ _1616_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xinput10 io_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_147_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3601_ mod.registers.r5\[4\] _0440_ _3292_ mod.registers.r11\[4\] _0571_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3348__A3 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _1547_ _1549_ _1550_ _1098_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6690__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6320_ _2759_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3532_ _3282_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6251_ _2888_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3463_ _3281_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ net12 _2142_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3505__B1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ mod.pc_1\[5\] _2869_ _2864_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3394_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _2005_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _2008_ _2009_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4835__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6470__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _0955_ _0561_ _0720_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _2424_ _2694_ _2698_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4233__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4917_ _1886_ _1883_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4784__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2655_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ mod.ldr_hzd\[13\] _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _1165_ _1485_ _1369_ _1185_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6518_ _3092_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _2715_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3914__I _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3511__A3 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6213__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4224__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__B2 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5972__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A1 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4160__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6906__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _2600_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _2531_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5963__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4702_ _1128_ _1669_ _1573_ _1330_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5682_ mod.registers.r8\[7\] _2510_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4633_ _1596_ _1601_ _1602_ _0917_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4518__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4564_ _1362_ _1533_ _0812_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5191__A2 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6303_ _2760_ _2959_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3515_ _3181_ _3197_ _3158_ _3184_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4495_ _1302_ _1464_ _1246_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout92_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6234_ mod.instr\[6\] _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3446_ _3285_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3377_ mod.instr_2\[2\] _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5116_ _2075_ _0958_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _2767_ _2799_ _2778_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _2010_ _1994_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4454__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6998_ _0096_ net218 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5949_ _2680_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5954__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__CLK net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__C2 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_303 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_314 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_325 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_336 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_347 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_358 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_369 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6198__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3708__B1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5173__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3300_ _3153_ _3154_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _3245_ _0896_ _0898_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6425__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _0019_ net202 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6852_ _0353_ net198 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6189__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _2566_ _2591_ _2595_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _0287_ net44 mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5936__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4334__B _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ mod.registers.r12\[15\] _0962_ _0964_ mod.registers.r15\[15\] _0965_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5734_ _2548_ _2541_ _2549_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _1572_ _1582_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6361__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _2445_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4547_ _1513_ _1516_ _1301_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4478_ _1445_ _1446_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6217_ mod.instr\[2\] _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ _3275_ _3277_ _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_89_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3478__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__B2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6148_ _2102_ _2824_ _2844_ _2789_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6416__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _1943_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5854__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3374__I _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6104__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4115__B1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4666__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout142_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ mod.registers.r13\[12\] _0745_ _0746_ mod.registers.r1\[12\] _0749_ _0750_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5450_ mod.registers.r3\[15\] _2350_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5381_ _2205_ _2309_ _2311_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4332_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout208 net212 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout219 net221 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4263_ _1113_ _0953_ _0957_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _2723_ mod.pc0\[0\] _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4194_ _3245_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4409__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _0405_ net152 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6835_ _0336_ net190 mod.pc0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5909__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6766_ _0270_ net60 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5385__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ _3250_ _0463_ _0919_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5717_ _2536_ _2530_ _2537_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6697_ _0201_ net111 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5674__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5648_ _2428_ _2486_ _2491_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5137__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5579_ _2386_ _2446_ _2449_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3320__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3871__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5376__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3926__A3 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4351__A3 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3311__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 io_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3862__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _1916_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6797__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3901_ mod.registers.r5\[9\] _0547_ _0548_ mod.registers.r7\[9\] _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4881_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6620_ _0124_ net134 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4024__C1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _3120_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3763_ _0503_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5502_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6482_ _3078_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6316__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3694_ mod.registers.r13\[3\] _0541_ _0542_ mod.registers.r1\[3\] _0663_ _0664_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5433_ _2331_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5364_ _2159_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__I _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4315_ _1182_ _1278_ _1282_ _1274_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _2163_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6258__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4246_ mod.registers.r8\[12\] _0968_ _0981_ mod.registers.r9\[12\] _1216_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _1144_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3853__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5055__B2 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _0322_ net40 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _0253_ net42 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A1 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5294__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4416__C _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3780__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout105_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3562__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4100_ _0688_ _0689_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _1135_ _0954_ _0957_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5285__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ mod.registers.r12\[14\] _0962_ _0996_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_84_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3835__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5037__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5489__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ _2708_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5588__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3599__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1797_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3599__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4260__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6537__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _3160_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3815_ mod.registers.r11\[14\] _0735_ _0746_ mod.registers.r1\[14\] _0785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6603_ _3149_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4795_ _1699_ _1764_ _1247_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4012__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ mod.registers.r15\[10\] _3107_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _3065_ _3067_ _3057_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3677_ _0609_ _0433_ _0417_ _0563_ _0610_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__6812__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ mod.registers.r3\[1\] _2332_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6396_ _0758_ _2953_ _3019_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5173__B _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4568__I _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ mod.registers.r1\[13\] _2277_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3472__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__A3 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ _2008_ _2210_ _2208_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6962__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ _1197_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4251__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3647__I _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4003__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4554__A3 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3514__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3817__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4490__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__C1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6835__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3600_ mod.registers.r12\[4\] _0437_ _0428_ mod.registers.r9\[4\] _0570_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput11 io_in[1] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _1547_ _0944_ _0938_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5742__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3531_ mod.registers.r8\[6\] _3272_ _0500_ mod.registers.r10\[6\] _0501_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__3753__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6250_ mod.instr\[10\] _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3462_ mod.registers.r9\[0\] _0428_ _0431_ mod.registers.r3\[0\] _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5201_ _1886_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3505__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3505__B2 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__B1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6181_ _1980_ _2868_ _2870_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3393_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _2056_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ mod.pc_2\[6\] _2009_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4014_ _0970_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4481__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ mod.registers.r14\[10\] _2695_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5430__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ mod.valid2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5896_ _2652_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ mod.ldr_hzd\[12\] _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4778_ _1384_ _1740_ _1742_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5733__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _2399_ _3093_ _3099_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3729_ _0695_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _3055_ _3044_ _3037_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5497__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6379_ _2713_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3511__A4 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5249__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3680__B1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6858__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5972__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5724__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A3 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__B1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4001__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4160__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4160__B2 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6129__S _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6452__A3 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5660__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout172_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5767__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4846__S0 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ _2529_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5963__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _1126_ _1371_ _1670_ _1186_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5681_ _2411_ _2509_ _2513_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4632_ _0901_ _1564_ _1566_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ _0828_ _0553_ _0773_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5191__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3514_ _0482_ _0483_ mod.registers.r13\[1\] _0477_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6302_ _1792_ _2958_ _2951_ mod.instr\[1\] _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4494_ _1224_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6233_ _2906_ _2901_ _2907_ _2905_ _2898_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3445_ _3284_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_143_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4151__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6164_ _2857_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout85_I net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3376_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ mod.pc_2\[10\] _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _2792_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3750__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ mod.pc_2\[5\] _1991_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5651__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _0095_ net220 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__A1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _2399_ _2681_ _2687_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5879_ mod.registers.r12\[10\] _2641_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A3 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4142__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__B2 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_304 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_315 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_326 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_337 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_348 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_359 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5642__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6680__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6192__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6198__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5587__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5945__A2 _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3708__A1 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3708__B2 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6211__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5881__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5633__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _0018_ net202 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _0352_ net198 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6189__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5802_ mod.registers.r10\[14\] _2592_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6782_ _0286_ net43 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5936__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3994_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3947__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ mod.registers.r9\[7\] _2542_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _2500_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4615_ _1300_ _1582_ _1584_ _3250_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5595_ _2414_ _2453_ _2458_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4350__B _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6361__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4546_ _1249_ _1515_ _1252_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ _0716_ _1310_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3428_ mod.instr_2\[13\] _3268_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6216_ _2893_ _2719_ _2894_ _2892_ _2855_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4675__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _2842_ _2843_ _2818_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3359_ mod.registers.r12\[0\] _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _2768_ _2004_ mod.pc\[2\] _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5029_ _1992_ _1975_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3650__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3655__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__B2 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4666__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__B _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3390__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__B1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5918__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3929__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3565__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4400_ _0932_ _0936_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4354__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ mod.registers.r2\[4\] _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4262_ _0779_ _0789_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout209 net210 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6001_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4657__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ _0953_ _1091_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3865__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A3 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3617__B1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _0404_ net154 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout48_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6116__I _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _0335_ net190 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A2 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6765_ _0269_ net57 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3977_ _0922_ _0928_ _0941_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5716_ mod.registers.r9\[2\] _2532_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _0200_ net91 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ mod.registers.r7\[11\] _2487_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ mod.registers.r6\[0\] _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _1496_ _1497_ _1383_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6098__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3320__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__I _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3385__I _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A2 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5836__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__I mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3698__I0 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3847__B1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_92_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3900_ mod.registers.r9\[9\] _0544_ _0545_ mod.registers.r3\[9\] _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4880_ _3255_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3831_ _0690_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4024__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4024__C2 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4575__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ mod.des.des_dout\[13\] net16 _3119_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3762_ _0502_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5501_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ mod.des.des_dout\[2\] net18 _3075_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3693_ _0660_ _0433_ _0661_ _0563_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6316__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4327__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _2329_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6600__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _2154_ _2157_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _0826_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5294_ _2201_ _2236_ _2237_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4245_ mod.registers.r6\[12\] _0966_ _0967_ mod.registers.r5\[12\] _1215_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _3266_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__I mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6817_ _0321_ net41 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5685__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6748_ _0252_ net120 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _0183_ net95 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4318__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3933__I _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__A2 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__B _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A3 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4004__I _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4939__I _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _0997_ _0998_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5285__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3296__A1 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4245__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ mod.pc0\[0\] _1892_ _1898_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3599__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__B _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4863_ _1817_ _1832_ _0478_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6537__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ net8 mod.des.des_dout\[36\] _3136_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3814_ _0780_ _0781_ _0782_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4794_ _1273_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6533_ _2421_ _3106_ _3109_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3745_ _3246_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _3055_ _1862_ _3066_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_146_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3676_ mod.registers.r9\[2\] _0544_ _0545_ mod.registers.r3\[2\] _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _2177_ _2330_ _2333_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6395_ mod.pc_1\[13\] _2720_ _3017_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5173__C _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4720__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4720__B2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _2221_ _2007_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4228_ mod.registers.r11\[13\] _0974_ _0972_ mod.registers.r10\[13\] mod.registers.r4\[13\]
+ _0971_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4159_ mod.registers.r12\[8\] _1110_ _0879_ mod.registers.r7\[8\] _1129_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5028__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4533__B _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4539__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__B2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5200__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6637__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3514__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__B1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__C2 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3838__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6214__I mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 io_in[2] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout215_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3530_ _3278_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3461_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5200_ net12 _1883_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4163__C1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3505__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6180_ mod.pc_1\[4\] _2869_ _2864_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3392_ _3238_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4702__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _1932_ _1775_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_151_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _1208_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6455__B2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ _0973_ _0976_ _0979_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _2421_ _2694_ _2697_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5430__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _1788_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3441__A1 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5895_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _1812_ _1813_ _1814_ _1815_ _1805_ _1808_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A1 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _1436_ _1746_ _1433_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6516_ mod.registers.r15\[3\] _3095_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3744__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3728_ mod.registers.r4\[3\] _0696_ _0697_ mod.registers.r1\[3\] _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3483__I _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _2966_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3659_ mod.registers.r8\[2\] _0531_ _0532_ mod.registers.r10\[2\] _0629_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5497__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _3007_ _3000_ _3008_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ mod.registers.r1\[11\] _2246_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6446__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5249__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3680__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3680__B2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5421__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3393__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3499__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__B2 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4160__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__A1 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__A1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout165_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__S1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _1549_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5680_ mod.registers.r8\[6\] _2510_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _1342_ _1598_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6952__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4562_ _0691_ _1334_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4399__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _2955_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3513_ _3217_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4493_ _1184_ _1190_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6232_ mod.des.des_dout\[5\] _2896_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3444_ mod.registers.r11\[0\] _3292_ _0413_ mod.registers.r2\[0\] _0414_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6163_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3375_ mod.funct3\[1\] _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _1743_ _1747_ _1756_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6094_ _1979_ _2797_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4348__B _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout78_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _1178_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5651__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4862__I _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6996_ _0094_ net210 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5403__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ mod.registers.r14\[3\] _2683_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5878_ _2554_ _2640_ _2643_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5167__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ mod.ins_ldr_3 mod.valid_out3 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5890__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_305 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_316 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_327 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_338 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_349 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6825__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6975__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5158__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3708__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4905__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4947__I _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5881__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5633__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__B1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__C2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6850_ _0351_ net192 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4615__C _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _2564_ _2591_ _2594_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _0285_ net43 mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3993_ _0485_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5732_ _2235_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5663_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _0912_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5594_ mod.registers.r6\[7\] _2454_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _1263_ _1268_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _1341_ _1054_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6215_ mod.des.des_dout\[1\] _2889_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3427_ mod.registers.r8\[0\] _3273_ _3279_ mod.registers.r10\[0\] _3280_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5321__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4124__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6848__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5872__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6146_ _2833_ _2838_ _2841_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__B2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6077_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _1971_ _1972_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input10_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6998__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _0077_ net101 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4060__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3936__I _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__B _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4115__A2 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4666__A3 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3874__B2 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5615__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7003__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4007__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4051__A1 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6222__I mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout128_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5000__B1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4354__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _0911_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _1003_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _2711_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3865__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ _0636_ _0952_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input2_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3865__B2 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3617__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3617__B2 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _0403_ net155 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _0334_ net175 mod.valid1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _0268_ net121 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4042__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3976_ _3241_ _0945_ _0463_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5715_ _2193_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5790__A1 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3396__A3 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _0199_ net95 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3756__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5646_ _2425_ _2486_ _2490_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5542__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5577_ _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6590__I0 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6670__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4528_ _1495_ _1496_ _1497_ _1432_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_104_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _1300_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ mod.pc\[8\] _2048_ _1894_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3320__A3 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6307__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__C _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4033__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5781__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3666__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3792__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6089__A2 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4497__I _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3847__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3847__B2 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3698__I1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6217__I mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4960__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3830_ _0579_ _0799_ _3262_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4024__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4024__B2 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5772__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3761_ mod.registers.r8\[12\] _0729_ _0730_ mod.registers.r10\[12\] _0731_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4575__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5500_ _2161_ _2356_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6693__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__B1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6480_ _3077_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3692_ mod.registers.r15\[3\] _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _2236_ _2337_ _2342_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5524__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4327__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5362_ _2270_ _2296_ _2297_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4313_ _1177_ _1179_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5293_ mod.registers.r1\[7\] _2206_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4244_ mod.registers.r3\[12\] _0959_ _0960_ mod.registers.r2\[12\] _0964_ mod.registers.r15\[12\]
+ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_102_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ _0633_ _0712_ _1044_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6252__A2 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4263__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _0320_ net63 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__C _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6747_ _0251_ net120 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5763__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4091__B _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _0455_ _0459_ _0452_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6678_ _0182_ net90 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5629_ _2472_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6563__I0 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4006__B2 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5506__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6909__CLK net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4955__I _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout195_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _2706_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4245__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__B2 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4931_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5786__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ _3213_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _3148_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3813_ mod.registers.r7\[14\] _0743_ _0729_ mod.registers.r8\[14\] mod.registers.r12\[14\]
+ _0766_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5745__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _1741_ _1745_ _1166_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6532_ mod.registers.r15\[9\] _3107_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3744_ _0595_ _0699_ _0710_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_9_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _2147_ _3025_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3675_ mod.registers.r5\[2\] _0547_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ mod.registers.r3\[0\] _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _2123_ _2953_ _3018_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5345_ mod.des.des_dout\[34\] _2213_ _2280_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4720__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5276_ _1786_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4227_ mod.registers.r12\[13\] _0962_ _0959_ mod.registers.r3\[13\] _0960_ mod.registers.r2\[13\]
+ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_75_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6473__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ mod.pc_2\[3\] _0778_ _1057_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__B1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3944__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3514__A3 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__D _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4475__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6216__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4227__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5975__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3738__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[3] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4950__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout110_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ _0429_ _0410_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout208_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__B1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__C2 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3391_ _3233_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5130_ _2072_ _2073_ _2088_ _3156_ _2089_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__B _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _1909_ _1720_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6881__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ mod.registers.r13\[15\] _0980_ _0981_ mod.registers.r9\[15\] _0982_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5963_ mod.registers.r14\[9\] _2695_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5966__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5894_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4845_ mod.ldr_hzd\[3\] _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _1741_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _2396_ _3093_ _3098_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3727_ _0466_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3744__A3 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4941__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _1826_ _3047_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3658_ mod.pc_2\[2\] _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_115_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6377_ mod.pc_1\[6\] _3001_ _3004_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3589_ mod.registers.r14\[4\] _3283_ _3287_ mod.registers.r6\[4\] _0559_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3901__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5328_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _2178_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6604__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6382__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__A2 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6050__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__A1 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3499__A2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4719__B _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout190 net193 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout158_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4620__B2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _1469_ _1599_ _0668_ _0924_ _0725_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4901__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ _1342_ _1527_ _1530_ _1419_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _2760_ _2957_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3512_ _3183_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4492_ _1436_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6231_ mod.instr\[5\] _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3443_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4687__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _2151_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A3 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3374_ _3226_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5113_ _1156_ _1160_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6093_ _2768_ _2769_ mod.pc\[4\] _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ mod.pc_2\[6\] _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3759__I _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6995_ _0093_ net211 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6135__I _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5179__C _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5946_ _2396_ _2681_ _2686_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5877_ mod.registers.r12\[9\] _2641_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4828_ _1191_ _0907_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5167__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3494__I _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _1538_ _1301_ _1537_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _3029_ _3041_ _3038_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3350__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A2 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5214__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_306 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_317 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_328 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_339 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3405__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5884__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5158__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6355__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6107__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__A1 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5330__A2 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3341__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__B2 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ mod.registers.r10\[13\] _2592_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6780_ _0284_ net134 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _0888_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _2546_ _2541_ _2547_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6830__D _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6346__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6346__B2 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _1071_ _1452_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5593_ _2411_ _2453_ _2457_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4544_ _1269_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4109__B1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3580__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1072_ _1063_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ mod.instr\[1\] _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout90_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3426_ _3278_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3332__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ _2833_ _2838_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _3209_ _3187_ _3206_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5034__I mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6076_ _2781_ _1913_ _1797_ _2770_ _2775_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5085__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5027_ mod.pc_2\[4\] _1972_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6978_ _0076_ net102 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _2430_ _2673_ _2675_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4541__C _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__I _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4899__A1 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3874__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5076__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6942__CLK net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3929__A3 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5000__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__C _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4260_ _1227_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ _1152_ _1156_ _1160_ _1143_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__3865__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5067__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__B _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3617__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6901_ _0402_ net155 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _0333_ net176 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _0267_ net136 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3975_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ _2534_ _2530_ _2535_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6319__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _0198_ net90 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ mod.registers.r7\[10\] _2487_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__CLK net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _2444_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5542__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__I1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4527_ _1492_ _1444_ _1456_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4458_ _1296_ _3242_ _1399_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6965__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3409_ _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4389_ _1356_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6128_ mod.pc\[9\] _2065_ _1894_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5058__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ _2764_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4552__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4033__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3792__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3792__B2 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__I1 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4344__I0 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3847__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3480__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4024__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5221__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3760_ _0500_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3783__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3783__B2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3691_ _0417_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ mod.registers.r3\[7\] _2338_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6988__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3806__B _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ mod.registers.r1\[15\] _2277_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _1279_ _1280_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5292_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4243_ _1209_ _1210_ _1211_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _0595_ _1131_ _1142_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5312__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout53_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _0319_ net62 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4015__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _0250_ net117 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3958_ _0925_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3774__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6677_ _0181_ net91 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3889_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _2400_ _2473_ _2479_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6563__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4574__I0 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ mod.registers.r5\[12\] _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5279__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__B _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5451__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3462__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4006__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__B1 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6554__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout188_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4930_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6660__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4861_ _1781_ _1191_ _0907_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_32_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6600_ net7 mod.des.des_dout\[35\] _3136_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3812_ mod.registers.r3\[14\] _0752_ _0736_ mod.registers.r2\[14\] _0782_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5745__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _1436_ _1760_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6531_ _2416_ _3106_ _3108_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3743_ _0615_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_146_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3674_ mod.registers.r7\[2\] _0548_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6462_ _1817_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5413_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6393_ mod.pc_1\[12\] _2720_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ _2166_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _2171_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _1192_ _1193_ _1194_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_68_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5681__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4157_ _1125_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _0657_ _0658_ _0659_ _0664_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_55_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3995__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3995__B2 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6729_ _0233_ net112 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6161__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3514__A4 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3683__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3435__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5975__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5727__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3738__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3738__B2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 io_in[4] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout103_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__B2 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3390_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4966__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3870__I _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _2021_ _2022_ _2023_ net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4011_ _0603_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5797__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _2416_ _2694_ _2696_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3977__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4913_ _1801_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _2161_ _2624_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ mod.ldr_hzd\[2\] _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6391__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _1188_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6514_ mod.registers.r15\[2\] _3095_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3726_ _0465_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _3052_ _3053_ _3046_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6143__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3657_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4154__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6376_ _2008_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3588_ mod.registers.r7\[4\] _0442_ _3273_ mod.registers.r8\[4\] _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3901__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3901__B2 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5327_ mod.des.des_dout\[32\] _2248_ _2264_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5654__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4209_ _3239_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _2140_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5406__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4209__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6134__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4145__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__C _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5645__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4448__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout180 net182 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout191 net193 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A3 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5410__I _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3959__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4620__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout220_I net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4560_ _0811_ _1528_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _0480_ _3256_ mod.registers.r14\[1\] _0477_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4491_ _1459_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3442_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6230_ _2903_ _2901_ _2904_ _2905_ _2898_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _2131_ _2824_ _2853_ _2854_ _2855_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3373_ mod.funct3\[2\] _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6092_ _1962_ _2766_ _2796_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5636__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1932_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4645__B _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5320__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _0092_ net211 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5945_ mod.registers.r14\[2\] _2683_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4611__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5876_ _2550_ _2640_ _2642_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _1389_ _1788_ _1791_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__6364__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3775__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4375__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4758_ _1724_ _1384_ _1725_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ _0675_ _0676_ _0677_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_107_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5990__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4689_ _0942_ _0914_ _0915_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6428_ _1858_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5875__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6100__B mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6359_ _2872_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3886__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_307 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_318 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_329 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6871__CLK net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4118__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout170_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ mod.registers.r3\[15\] _0959_ _0960_ mod.registers.r2\[15\] _0961_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5730_ mod.registers.r9\[6\] _2542_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ _2357_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _1580_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5592_ mod.registers.r6\[6\] _2454_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ _1512_ _1439_ _1438_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4109__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__B2 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _1437_ _1256_ _1441_ _1443_ _1257_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5857__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6213_ _2887_ _2719_ _2890_ _2892_ _2855_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3425_ _3267_ _3269_ _3275_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6144_ _2101_ _2840_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3356_ _3158_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout83_I net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ mod.pc\[1\] _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5026_ _1163_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6744__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _0075_ net45 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6894__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ mod.registers.r13\[12\] _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__B _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ mod.registers.r12\[2\] _2629_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4348__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5848__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3859__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4520__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__A2 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__B1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6005__B _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4511__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ _1157_ _1158_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6767__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6900_ _0401_ net166 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4814__B3 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6831_ _0002_ _0006_ net217 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__4027__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6762_ _0266_ net136 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3974_ _0942_ _0943_ _0915_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4042__A3 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5713_ mod.registers.r9\[1\] _2532_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3539__B _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ _0197_ net91 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5644_ _2422_ _2486_ _2489_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4526_ _1259_ _1271_ _1151_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4750__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _1418_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5045__I _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4502__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3408_ _3253_ _3180_ _3222_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4388_ _1357_ _0840_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ _2817_ _2820_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ mod.registers.r6\[0\] _3186_ _3189_ mod.registers.r5\[0\] mod.registers.r2\[0\]
+ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6058_ _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _1953_ _1973_ _1954_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4833__B _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__A2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3792__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4344__I1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6246__B2 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4009__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3480__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__B _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3480__B2 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5221__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout133_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ mod.registers.r12\[3\] _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__I mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _0874_ _1121_ _1123_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5291_ mod.des.des_dout\[28\] _2188_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5288__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4242_ mod.registers.r12\[12\] _0962_ _0975_ mod.registers.r1\[12\] _1212_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _1021_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4637__C _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4799__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout46_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _0318_ net58 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _0249_ net121 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ _0926_ _0774_ _0453_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3774__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _0180_ net48 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3888_ _0843_ _3239_ _0852_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5627_ mod.registers.r7\[3\] _2475_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4184__C1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _2390_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4574__I1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4509_ _1329_ _1472_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ _2361_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4239__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4119__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5451__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3462__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4563__B _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3462__B2 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4962__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4714__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5413__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__A2 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6805__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ _1803_ _1811_ _1829_ _3244_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3811_ mod.registers.r15\[14\] _0765_ _0751_ mod.registers.r9\[14\] _0781_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6955__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _1273_ _1278_ _1759_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6530_ mod.registers.r15\[8\] _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3742_ mod.funct7\[0\] _0711_ _0617_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4699__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6461_ _3032_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3673_ _0629_ _0630_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5412_ _2328_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4705__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6392_ _2752_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ _2042_ _2241_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6458__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _2201_ _2218_ _2219_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5130__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4225_ mod.registers.r1\[13\] _0975_ _0981_ mod.registers.r9\[13\] _1195_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5130__B2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5681__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ _0873_ _1124_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_110_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ _0652_ _0653_ _0654_ _0655_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3778__I mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__B _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3444__B2 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4989_ _1952_ _1955_ _1794_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ _0232_ net93 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6659_ _0163_ net80 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6103__B _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4558__B _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3683__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3683__B2 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5424__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__B2 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3738__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4935__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 io_in[5] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4163__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__I mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4010_ _0608_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3674__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5961_ mod.registers.r14\[8\] _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4912_ _1830_ _1876_ _1881_ _1817_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _2568_ _2646_ _2651_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5179__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5179__B2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4843_ mod.ldr_hzd\[1\] _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4774_ _1102_ _1105_ _1279_ _1492_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6513_ _2393_ _3093_ _3097_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3725_ mod.registers.r3\[3\] _0694_ _0596_ mod.registers.r7\[3\] _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _2967_ _3041_ _3037_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3656_ _0625_ _0622_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5351__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _0580_ _3000_ _3006_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3587_ _0459_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5326_ _2166_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3901__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5257_ mod.des.des_dout\[25\] _2167_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4208_ _0424_ _0953_ _0956_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4892__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _1107_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5406__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4090__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5342__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5893__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4288__B _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__I _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5645__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout170 net173 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3656__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout181 net182 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout192 net193 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3408__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__B1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3959__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5581__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout213_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3510_ _3209_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4490_ _1224_ _1276_ _1286_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3441_ _3275_ _3277_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5333__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _2788_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3372_ _3154_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A1 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__B2 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5111_ _0000_ mod.des.des_counter\[1\] _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6091_ _0003_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5636__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _1685_ _1696_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__C _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _0091_ net213 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _2393_ _2681_ _2685_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ mod.registers.r12\[8\] _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6432__I _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4826_ _1794_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5572__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _1699_ _1723_ _1726_ _1247_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ mod.registers.r9\[1\] _0511_ _0500_ mod.registers.r10\[1\] _0678_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _1383_ _1650_ _1653_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6427_ _1814_ _3033_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3639_ mod.registers.r12\[2\] _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6358_ _2952_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3886__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5309_ _1972_ _2241_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3350__A3 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6289_ mod.des.des_dout\[20\] _2900_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_308 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_319 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5511__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6342__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5563__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4366__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3326__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5866__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3877__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6291__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout163_I net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _0701_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__B _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _2146_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _1267_ _1264_ _1266_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5554__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5591_ _2408_ _2453_ _2456_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _1448_ _1453_ _1454_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__A2 _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _1097_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ _2891_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3424_ _3276_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ mod.pc\[11\] _1914_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3355_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3332__A3 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6074_ _2765_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout76_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5025_ _1082_ _1087_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6034__A2 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _0074_ net41 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5793__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ _2655_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6162__I _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _2534_ _2627_ _2631_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5545__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4348__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _1390_ _1394_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5789_ _2550_ _2585_ _2587_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3859__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__B2 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6337__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__A1 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__B2 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5784__A1 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5536__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__A2 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6830_ _0001_ _0005_ net219 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__4027__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4027__B2 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5775__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _0265_ net121 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3973_ _0935_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5712_ _2185_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4042__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6692_ _0196_ net47 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5527__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ mod.registers.r7\[9\] _2487_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4525_ _0912_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4456_ _1235_ _1371_ _1424_ _1331_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3407_ _3254_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4502__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4387_ _0460_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ mod.pc\[9\] _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3710__B1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4386__B _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4266__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6861__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ mod.pc_2\[3\] _1951_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4018__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4833__C _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _0057_ net213 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5518__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5236__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__A2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4140__I _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__B1 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6067__I _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__A1 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__B2 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3480__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5509__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4980__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout126_I net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4310_ _0859_ _1144_ _1146_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5290_ _2231_ _2232_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ mod.registers.r14\[12\] _0977_ _0978_ mod.registers.r7\[12\] _1211_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__A1 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4172_ _1132_ _1133_ _1140_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4799__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5748__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _0317_ net62 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout39_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _0248_ net107 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3956_ _3246_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ _0179_ net47 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3887_ _0853_ _0854_ _0855_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5626_ _2397_ _2473_ _2478_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4184__B1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5920__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _2388_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4184__C2 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4508_ _1473_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _2359_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4439_ _0757_ _0774_ _1291_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _2808_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4239__B2 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3462__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5739__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A2 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4411__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__CLK net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3922__B1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3642__C _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5978__A1 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3453__A2 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3810_ mod.registers.r5\[14\] _0741_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4790_ _1278_ _1759_ _1273_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3741_ _3215_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _2716_ _3063_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3672_ _0498_ _0635_ _0639_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5411_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _2095_ _2953_ _3016_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5902__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3913__B1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5342_ _0758_ _2181_ _2214_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_154_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4929__B _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__B _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ mod.registers.r1\[5\] _2206_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4224_ mod.registers.r14\[13\] _0977_ _0889_ mod.registers.r13\[13\] _0978_ mod.registers.r7\[13\]
+ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5130__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _0873_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3444__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _1953_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6727_ _0231_ net97 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3939_ mod.funct7\[1\] _0905_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6658_ _0162_ net76 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _2431_ _2465_ _2467_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _3135_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__A3 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3683__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4632__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6137__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 io_in[6] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3371__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout193_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3674__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6922__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6255__I mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _2682_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _1877_ _1878_ _1879_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5891_ mod.registers.r12\[15\] _2647_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5179__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ mod.ldr_hzd\[0\] _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4773_ _1740_ _1742_ _1699_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6604__RN _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4503__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ mod.registers.r15\[1\] _3095_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3724_ _0471_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _0495_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6443_ _1822_ _3047_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6374_ mod.pc_1\[5\] _3001_ _3004_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3586_ _0455_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4659__B _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ _2009_ _2241_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5256_ _2181_ _1968_ _2173_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6300__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _1152_ _1171_ _1176_ _1143_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5187_ net11 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3665__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ mod.registers.r3\[9\] _0694_ _0882_ mod.registers.r5\[9\] _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3789__I _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6165__I _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input19_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4069_ mod.registers.r1\[6\] _0466_ _3204_ mod.registers.r8\[6\] _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3417__A2 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4614__A1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4090__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4413__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A3 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3353__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6945__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout160 net168 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout171 net173 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4853__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout182 net183 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout193 net194 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3699__I mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6075__I mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3408__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__B2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__A3 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3813__C1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5581__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__A3 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3440_ _3284_ _3268_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6530__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3371_ _3180_ _3222_ _3223_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _1908_ _2055_ _2069_ _0001_ _2070_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ _2792_ _2794_ _2773_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5097__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5041_ _1916_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3402__I mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ _0090_ net214 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ mod.registers.r14\[1\] _2683_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4434__S _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5874_ _2628_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__B2 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ mod.pc_2\[0\] _1078_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5021__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6818__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5572__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _1724_ _1725_ _1302_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3707_ mod.registers.r5\[1\] _0517_ _0518_ mod.registers.r7\[1\] _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _1243_ _1655_ _1656_ _1433_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3638_ _3210_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6426_ _3035_ _3039_ _3023_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6521__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6968__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3335__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3569_ _0533_ _0536_ _0537_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_88_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _2992_ _2994_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3886__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5308_ _2191_ _2055_ _2209_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6288_ mod.instr\[20\] _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_309 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5239_ _2165_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__I _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__I1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4344__S _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5012__A1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4143__I _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5563__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6512__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5315__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4299__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__B2 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3877__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3341__A4 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4826__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6291__A3 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout156_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5149__I _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _1449_ _1451_ _1452_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5590_ mod.registers.r6\[5\] _2454_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5554__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4541_ _1494_ _1498_ _1499_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4762__B1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3892__I mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4472_ _1048_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6211_ net13 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3423_ mod.instr_2\[10\] _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6142_ _2832_ _2839_ _2831_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3354_ _3183_ _3184_ _3206_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3332__A4 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6073_ _2774_ _2777_ _2779_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1987_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout69_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _0073_ net41 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4672__B _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5926_ _2653_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5857_ mod.registers.r12\[1\] _2629_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4808_ _1376_ _1698_ _1758_ _1775_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5788_ mod.registers.r10\[8\] _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4739_ _1635_ _1636_ _1343_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6409_ _1850_ _2883_ _3027_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5522__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4808__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6554__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__B _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5784__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6528__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5472__A1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4275__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6663__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6263__I mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6760_ _0264_ net102 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _3248_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5711_ _2527_ _2530_ _2533_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6691_ _0195_ net47 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5642_ _2417_ _2486_ _2488_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _2299_ _2356_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5607__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _1491_ _1493_ _1242_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4455_ _1004_ _0934_ _1246_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3406_ _3255_ _3256_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4386_ _0813_ _0814_ _0826_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3710__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6125_ _2818_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3337_ _3182_ _3159_ _3163_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3710__B2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6056_ _2725_ _1899_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4266__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ mod.pc_2\[3\] _1951_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A2 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6958_ _0056_ net215 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5909_ _2402_ _2661_ _2663_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6889_ _0390_ net171 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4726__B1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4421__I _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3701__A1 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6348__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3701__B2 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4257__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4009__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5206__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__S _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4331__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3940__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ mod.registers.r11\[12\] _0974_ _0980_ mod.registers.r13\[12\] _1210_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5693__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4171_ mod.registers.r2\[8\] _0893_ _0468_ mod.registers.r5\[8\] mod.registers.r11\[8\]
+ _0605_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_110_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5445__A1 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _0316_ net122 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5748__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6743_ _0247_ net108 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3955_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6674_ _0178_ net40 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3886_ mod.registers.r5\[8\] _0440_ _0413_ mod.registers.r2\[8\] _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5625_ mod.registers.r7\[2\] _2475_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5337__I _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4184__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4184__B2 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5556_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5920__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4507_ _0811_ _1474_ _1475_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5487_ _2268_ _2373_ _2378_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4438_ _1404_ _1407_ _1351_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4369_ _1336_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6108_ _2016_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _2139_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3521__S _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5021__B _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5739__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4411__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A2 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3922__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3922__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3990__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5978__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6701__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__B _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4402__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _0702_ _0704_ _0707_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_13_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__I mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ _0637_ _0445_ mod.registers.r2\[2\] _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6851__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6390_ mod.pc_1\[11\] _2720_ _3012_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3913__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3913__B2 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _2182_ _2122_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4469__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ mod.registers.r6\[13\] _0966_ _0967_ mod.registers.r5\[13\] _1193_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3677__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ _1121_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__A1 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4437__S _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4085_ _0759_ _0620_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5620__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6091__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4680__B _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _1051_ _1935_ _1917_ _1937_ _1938_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6394__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6451__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6726_ _0230_ net92 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3601__B1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3938_ _0902_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6657_ _0161_ net85 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3869_ mod.pc_2\[10\] _0778_ _0833_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ mod.registers.r6\[12\] _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6588_ _3141_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5539_ _2388_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__I _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6724__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 io_in[7] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6137__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3371__A2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5648__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3659__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout186_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__B1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ _1815_ _1814_ _1813_ _1812_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_45_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ _2566_ _2646_ _2650_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _1804_ _1806_ _0661_ _1807_ _1809_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__6271__I mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ _1741_ _1281_ _1650_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6511_ _2385_ _3093_ _3096_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3723_ _0627_ _0668_ _0686_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6442_ _3050_ _3051_ _3046_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3654_ _0497_ _0555_ _0594_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5887__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _3003_ _3000_ _3005_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3898__B1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3585_ _0526_ _0527_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ _2191_ _2090_ _2214_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout99_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5255_ _1971_ _2182_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4206_ _1172_ _1173_ _1174_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_87_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5186_ _2138_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3665__A3 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ mod.registers.r10\[9\] _1106_ _0703_ mod.registers.r9\[9\] _1107_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ mod.registers.r3\[6\] _0471_ _0465_ mod.registers.r4\[6\] _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5811__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6897__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__B1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _0213_ net91 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6119__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5525__I _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A4 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3353__A2 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout150 net158 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout161 net168 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout172 net174 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout183 net184 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout194 net201 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6055__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4066__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__A1 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3408__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__B1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3813__C2 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6602__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A3 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5869__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout101_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3370_ _3153_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _1787_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__B _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__I mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6046__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6991_ _0089_ net214 mod.des.des_dout\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _2385_ _2681_ _2684_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ _2626_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6349__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4514__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _1792_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5021__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _1204_ _1459_ _1292_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3706_ mod.registers.r14\[1\] _0502_ _3291_ mod.registers.r11\[1\] _0676_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4780__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ _1506_ _1493_ _1651_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6425_ _3029_ _3036_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3637_ _3207_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6356_ _0955_ _2989_ _2962_ mod.instr\[20\] _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3568_ mod.registers.r4\[7\] _0508_ _3237_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ mod.pc_2\[9\] _2221_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6287_ _2946_ _2889_ _2947_ _2941_ _2742_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3499_ mod.registers.r2\[1\] _3191_ _0468_ mod.registers.r5\[1\] _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _2164_ _2186_ _2187_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _2124_ _2111_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6037__A1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4424__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3877__A3 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__B1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _1504_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4471_ _1438_ _1439_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6210_ mod.des.des_dout\[0\] _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3422_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6141_ _2834_ _2836_ _2838_ _2817_ _2773_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3353_ _3161_ mod.instr_2\[16\] _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6072_ mod.pc\[1\] _2774_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5114__B _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _3243_ _1554_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3413__I _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6019__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4445__S _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6974_ _0072_ net45 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5925_ _2427_ _2667_ _2672_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _2527_ _2627_ _2630_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4807_ _1392_ _1395_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5787_ _2573_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4202__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ _1429_ _0901_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _0717_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ mod.rd_3\[0\] _2884_ _3017_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4505__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _2978_ _2983_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6258__B2 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4419__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3323__I mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__B _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3993__I _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__C _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__B2 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6808__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5472__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6421__A1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6958__CLK net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3971_ _0929_ _0934_ _0685_ _0938_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ mod.registers.r9\[0\] _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6690_ _0194_ net40 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5641_ mod.registers.r7\[8\] _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5572_ _2442_ _2432_ _2443_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ _1102_ _1105_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4454_ _1420_ _1421_ _1423_ _1340_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__A1 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3405_ mod.funct3\[2\] _3232_ _3257_ _3234_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_131_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4385_ _1353_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6124_ _2050_ _2780_ _2823_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout81_I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3336_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3710__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6055_ _2734_ _2134_ _2763_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _1122_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _0055_ net219 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ mod.registers.r13\[4\] _2662_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6888_ _0389_ net171 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5839_ _2598_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4726__A1 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__B2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5533__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__S _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__B _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__B1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__A1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5142__A1 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6539__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6630__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _1134_ _1137_ _1138_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6780__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _0315_ net120 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6742_ _0246_ net103 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3954_ _0923_ _0808_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6673_ _0177_ net48 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5618__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3885_ mod.registers.r14\[8\] _3283_ _0428_ mod.registers.r9\[8\] _0855_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _2394_ _2473_ _2477_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4708__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5555_ _2275_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4184__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5381__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _1316_ _0927_ _1350_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ mod.registers.r4\[11\] _2374_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6449__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _1405_ _0462_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5353__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4368_ _1337_ _0724_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _2802_ _1885_ mod.pc\[6\] _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3319_ _3158_ _3159_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0899_ _1251_ _1075_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6038_ _2730_ _2053_ _2751_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6184__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5021__C _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A4 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4860__C _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6133__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3922__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5263__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3686__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5427__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3453__A4 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3670_ _0631_ _0562_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ _2270_ _2276_ _2278_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3913__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ mod.des.des_dout\[26\] _2188_ _2212_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4222_ mod.registers.r15\[13\] _0964_ _0968_ mod.registers.r8\[13\] _1192_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3677__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3677__B2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ _0577_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3429__A1 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4084_ _1051_ _0499_ _1052_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_110_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_290 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout44_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _1051_ _1935_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6725_ _0229_ net92 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3937_ _0904_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3601__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3601__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _0160_ net128 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3868_ _0834_ _0835_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_149_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _2447_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5354__A1 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ net19 mod.des.des_dout\[29\] _3137_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3799_ mod.registers.r9\[13\] _0428_ _0752_ mod.registers.r3\[13\] _0769_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5538_ _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6179__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _2361_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5657__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3668__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3331__I mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5593__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5258__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 io_in[8] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5345__A1 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5648__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3659__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__B2 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__B1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4337__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__B2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4781__B _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6699__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4840_ mod.ldr_hzd\[10\] _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5584__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _1272_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ mod.registers.r15\[0\] _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3595__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3722_ _0691_ _0622_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _2967_ _3036_ _3037_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5336__A1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3653_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3347__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ mod.pc_1\[4\] _3001_ _3004_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3584_ _0529_ _0551_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3898__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3898__B2 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5323_ mod.pc_2\[11\] _2169_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5254_ _2163_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4205_ mod.registers.r12\[11\] _1110_ _0882_ mod.registers.r5\[11\] _0696_ mod.registers.r4\[11\]
+ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_69_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ _1781_ net31 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _3195_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3665__A4 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _1034_ _1035_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4075__A1 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__B2 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _0954_ _0492_ _1936_ _0669_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_6708_ _0212_ net50 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5327__A1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6639_ _0143_ net84 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_94_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout151 net153 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout162 net167 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout173 net174 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout184 net185 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout195 net197 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6841__CLK net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__B2 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3996__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3813__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__B2 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6602__I1 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6483__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4057__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _0088_ net213 mod.des.des_dout\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5941_ mod.registers.r14\[0\] _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__I mod.instr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5872_ _2548_ _2634_ _2639_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _0903_ _0906_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4754_ _1287_ _1293_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_159_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3705_ mod.registers.r15\[1\] _0514_ _0512_ mod.registers.r3\[1\] _0675_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5309__A1 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ _1651_ _1506_ _1493_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4780__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3636_ mod.registers.r11\[2\] _0605_ _0473_ mod.registers.r8\[2\] _0606_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6424_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _2992_ _2993_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3335__A3 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3567_ mod.registers.r11\[7\] _0505_ _0506_ mod.registers.r2\[7\] _0537_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5306_ _2165_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ mod.des.des_dout\[19\] _2900_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3498_ _3188_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5237_ mod.registers.r1\[1\] _2179_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4296__B2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _2123_ _1089_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ mod.funct7\[2\] _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ mod.pc_2\[9\] _1233_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6596__I0 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4220__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6568__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__A4 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__I _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4287__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4039__B2 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6587__I0 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4211__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4762__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout211_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _1253_ _1099_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ mod.instr_2\[11\] _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3352_ mod.registers.r11\[0\] _3202_ _3204_ mod.registers.r8\[0\] _3205_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6277__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6071_ _2753_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5022_ _3154_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6973_ _0071_ net59 mod.registers.r15\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5924_ mod.registers.r13\[11\] _2668_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5855_ mod.registers.r12\[0\] _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _1394_ _1698_ _1758_ _1775_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4202__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _2571_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4202__B2 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4737_ _1701_ _1702_ _1384_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4753__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _0811_ _1635_ _1636_ _1637_ _1468_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3619_ mod.registers.r13\[5\] _0446_ _0448_ mod.registers.r1\[5\] _0589_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4505__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _3025_ _3026_ _3023_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _0809_ _1532_ _1534_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_134_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6338_ _0846_ _2982_ _2979_ mod.instr\[13\] _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6258__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _2741_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A3 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3492__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4441__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5941__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4103__C _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6249__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__I _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout161_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4432__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4983__A2 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5640_ _2474_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5571_ mod.registers.r5\[15\] _2433_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5932__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3943__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4522_ _1490_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4453_ _1242_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4948__C _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3404_ mod.instr_2\[2\] mod.instr_2\[0\] _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4384_ _0683_ _0684_ _0859_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6123_ _2765_ _2821_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3335_ _3166_ _3167_ _3175_ _3187_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6054_ mod.pc0\[13\] _2723_ _2754_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5999__A1 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ mod.pc_2\[4\] _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6902__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6956_ _0054_ net148 mod.ldr_hzd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _2655_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4974__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6887_ _0388_ net171 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3631__C1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6176__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ _2558_ _2612_ _2617_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4187__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _2527_ _2572_ _2575_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5151__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__B _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5454__A3 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__B2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__A2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__I _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6581__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__A2 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6380__I _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5914__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4717__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6925__CLK net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6810_ _0314_ net117 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4405__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6741_ _0245_ net107 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ _0625_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _0176_ net53 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3884_ mod.registers.r13\[8\] _0447_ _3279_ mod.registers.r10\[8\] _0854_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5905__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5623_ mod.registers.r7\[1\] _2475_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4708__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3419__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5554_ _2428_ _2418_ _2429_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5381__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4505_ _1401_ _1310_ _0575_ _0812_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5485_ _2261_ _2373_ _2377_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _0801_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4367_ _1250_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6106_ _2783_ _2791_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3318_ mod.registers.r3\[0\] _3165_ _3170_ mod.registers.r7\[0\] _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4298_ _1264_ _1266_ _1267_ _1260_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _2729_ mod.pc0\[8\] _2731_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4644__B2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_162_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6939_ _0037_ net162 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6149__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3329__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4869__B _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5544__I _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6576__S _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3686__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__A1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _2213_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ _0720_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6486__S _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3677__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _0637_ _0897_ _1044_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6076__B1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6285__I mod.instr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4083_ _0644_ _0645_ _0646_ _0648_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_83_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_280 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_291 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _0651_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6724_ _0228_ net49 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3936_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3601__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _0159_ net159 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3867_ mod.registers.r13\[10\] _0745_ _0746_ mod.registers.r1\[10\] _0837_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5606_ _2445_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5354__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6586_ _3140_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3798_ mod.registers.r13\[13\] _0447_ _0449_ mod.registers.r1\[13\] _0768_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3365__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5537_ _2244_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5106__A2 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6303__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _2359_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5399_ _2303_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3668__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4865__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6620__CLK net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5593__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput19 io_in[9] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3522__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4608__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__C1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4770_ _1738_ _1739_ _1167_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5584__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3595__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6440_ _1824_ _3047_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3652_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5336__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3347__A1 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3347__B2 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6371_ _2872_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5184__I _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3583_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3898__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5322_ _2238_ _2261_ _2262_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _2164_ _2199_ _2200_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4204_ mod.registers.r8\[11\] _0706_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5184_ _2137_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__A3 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4135_ _1031_ _0525_ _1103_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_95_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ mod.registers.r5\[6\] _3189_ _3199_ mod.registers.r9\[6\] _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6643__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4968_ _3229_ _0954_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ _0211_ net49 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _3211_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4899_ _1861_ _1867_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6524__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6638_ _0142_ net87 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5327__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3607__I _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _3130_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout130 net131 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout141 net142 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout152 net157 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout163 net167 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout174 net184 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout185 net203 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3342__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout196 net197 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4066__A2 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6515__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5732__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout191_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6666__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5871_ mod.registers.r12\[7\] _2635_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _1191_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3568__A1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__B1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4753_ _1722_ _1204_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5907__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3704_ _0670_ _0671_ _0672_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4684_ _1650_ _1653_ _1429_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6423_ mod.instr_2\[6\] _3025_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3635_ _3201_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6354_ mod.funct7\[1\] _2989_ _2962_ mod.instr\[19\] _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ mod.registers.r14\[7\] _0534_ _0535_ mod.registers.r6\[7\] _0536_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3335__A4 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3871__B _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _2238_ _2245_ _2247_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ mod.instr\[19\] _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3497_ mod.registers.r4\[1\] _0465_ _0466_ mod.registers.r1\[1\] _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5236_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4258__I _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _2123_ _1089_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _1082_ _1087_ _0457_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5098_ _2057_ _2045_ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ mod.registers.r14\[7\] _0607_ _0596_ mod.registers.r7\[7\] _1019_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4599__A3 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__C1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6596__I1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__S0 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6141__C _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5181__B1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__I _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6689__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5484__A1 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4287__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4039__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3798__B2 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6587__I1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4211__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6558__I _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6070_ _2771_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ _1908_ _1968_ _1984_ _1986_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _0070_ net59 mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5778__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__C _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5923_ _2424_ _2667_ _2671_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ _2628_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _1762_ _1765_ _1766_ _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5785_ _2548_ _2579_ _2584_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4202__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4736_ _1699_ _1701_ _1702_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ _1350_ _1334_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__CLK net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ mod.ins_ldr_3 _2995_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3618_ mod.registers.r5\[5\] _0439_ _0441_ mod.registers.r7\[5\] _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5702__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__B _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4598_ _1524_ _1526_ _0623_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6337_ _2860_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3549_ mod.registers.r5\[6\] _0517_ _0518_ mod.registers.r7\[6\] _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_88_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6268_ mod.des.des_dout\[14\] _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6981__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5466__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4269__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _2169_ _1387_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4808__A4 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ mod.pc_1\[11\] _2877_ _2880_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A3 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A2 _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__A2 _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__B1 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3468__B1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3530__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4432__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout154_I net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6854__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2441_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5932__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3943__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _1102_ _1105_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3943__B2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4452_ _0923_ _1305_ _0950_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5696__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__I mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _3187_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _0926_ _0774_ _0874_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5192__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6122_ _2753_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _3176_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6053_ _2760_ _2762_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _1794_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout67_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4536__I _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6955_ _0053_ net147 mod.ldr_hzd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5906_ _2653_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6886_ _0387_ net170 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3631__B1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3631__C2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ mod.registers.r11\[11\] _2613_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6176__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5367__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4187__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4187__B2 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ mod.registers.r10\[0\] _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1307_ _1598_ _1688_ _1328_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5699_ _2436_ _2521_ _2524_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5687__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5439__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A2 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__C _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__B2 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6727__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5678__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4130__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3689__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5602__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _0244_ net68 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3952_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3613__B1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6671_ _0175_ net53 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6158__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3883_ mod.registers.r1\[8\] _0449_ _0431_ mod.registers.r3\[8\] _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4169__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _2386_ _2473_ _2476_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ mod.registers.r5\[11\] _2419_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _0461_ _1054_ _0682_ _0923_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5484_ mod.registers.r4\[10\] _2374_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5669__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _0461_ _1054_ _0682_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4366_ _0878_ _1241_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6105_ _1979_ _2797_ _1998_ _2803_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3317_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5650__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _1055_ _1061_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6094__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6036_ _2743_ _2750_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _0036_ net163 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _0370_ net188 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3907__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3686__A3 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5832__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6388__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5060__A2 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5735__I _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4571__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4323__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4220_ _1180_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4795__B _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3677__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4151_ _3253_ _1109_ _1120_ _1021_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__6076__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _0629_ _0630_ _0642_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_95_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5823__A1 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3429__A3 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_270 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_281 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_292 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _1145_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6723_ _0227_ net39 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3935_ _3231_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _0158_ net160 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3866_ mod.registers.r5\[10\] _0741_ _0743_ mod.registers.r7\[10\] _0836_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5605_ _2428_ _2459_ _2464_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6585_ net18 mod.des.des_dout\[28\] _3137_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3797_ mod.registers.r15\[13\] _0765_ _0766_ mod.registers.r12\[13\] _0767_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5536_ _2414_ _2404_ _2415_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5467_ _2199_ _2360_ _2366_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ mod.valid2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5398_ _2301_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4865__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _1074_ _0527_ _0573_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5814__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _2734_ mod.pc0\[3\] _2737_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3825__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__I _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3803__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4069__B1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5805__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__B1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3816__C2 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3678__C _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6230__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _0688_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3595__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _0578_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6533__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3347__A2 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1971_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3582_ _3261_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ mod.registers.r1\[10\] _2246_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6497__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ mod.registers.r1\[3\] _2179_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4203_ mod.registers.r15\[11\] _0884_ _1106_ mod.registers.r10\[11\] _1173_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3713__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _1792_ _0907_ _1887_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _1030_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ mod.registers.r15\[6\] _0963_ _3186_ mod.registers.r6\[6\] _1035_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4544__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6221__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6938__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4967_ _1025_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6706_ _0210_ net39 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3918_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4898_ mod.ldr_hzd\[14\] _1857_ _1853_ mod.ldr_hzd\[13\] mod.ldr_hzd\[12\] _1856_
+ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6637_ _0141_ net84 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3849_ _0815_ _0816_ _0817_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_164_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4535__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ mod.des.des_dout\[21\] net6 _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _2204_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6499_ mod.des.des_dout\[10\] net8 _3085_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5324__B _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout120 net123 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3623__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout142 net143 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout153 net157 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout164 net166 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout175 net176 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout186 net189 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout197 net200 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4390__S _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4526__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3533__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout184_I net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _2546_ _2634_ _2638_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4821_ _1790_ _1387_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3568__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4765__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4752_ _1222_ _1463_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4765__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ mod.registers.r4\[1\] _0419_ _3264_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _1651_ _1280_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6422_ _1854_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4517__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3634_ mod.registers.r10\[2\] _0602_ _0603_ mod.registers.r9\[2\] _0604_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4517__B2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6353_ _2707_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3565_ _3286_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ mod.registers.r1\[8\] _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6284_ _2944_ _2937_ _2945_ _2941_ _2742_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_fanout97_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3496_ _3177_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ mod.des.des_dout\[22\] _2167_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3443__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6610__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _0727_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4117_ _1083_ _1084_ _1085_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5097_ mod.pc_2\[8\] _2042_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4048_ _1011_ _1012_ _1016_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__B1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _2719_ _2721_ _2716_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__C2 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4756__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__S1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4508__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5181__B2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6433__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3798__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A3 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5743__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__C _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3350_ _3196_ _3197_ _3172_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4359__I _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5020_ _0886_ _0895_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6783__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _0069_ net60 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5922_ mod.registers.r13\[10\] _2668_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4986__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5853_ _2625_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4738__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4804_ _1659_ _1767_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4822__I _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5784_ mod.registers.r10\[7\] _2580_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6242__C _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _1437_ _1703_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3438__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _0802_ _1356_ _1364_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _1831_ _2856_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3617_ mod.registers.r9\[5\] _0427_ _0430_ mod.registers.r3\[5\] _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5163__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _0901_ _1565_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6336_ _2978_ _2981_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4910__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3548_ _0441_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _2717_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5466__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _1786_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6198_ _2085_ _2876_ _2881_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ _1932_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__CLK net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5154__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3704__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__A1 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__B2 mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4968__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout147_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5393__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _1148_ _1149_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3943__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _0924_ _0790_ _0800_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_144_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5696__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3402_ mod.instr_2\[3\] _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4382_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6121_ _2816_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6052_ _2746_ mod.pc0\[12\] _2761_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _3155_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3721__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4959__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _0052_ net148 mod.ldr_hzd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5905_ _2399_ _2654_ _2660_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3631__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6885_ _0386_ net163 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__B2 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6679__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3596__C _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5836_ _2556_ _2612_ _2616_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4187__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5384__A1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4718_ _1343_ _1686_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5698_ mod.registers.r8\[13\] _2522_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ _1514_ _0945_ _1366_ _1477_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5687__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _2961_ _2970_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4111__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5611__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5558__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3622__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__I _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5127__B2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3689__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3689__B2 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3742__S _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3541__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__B2 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6821__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _0724_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_16_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3613__A1 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3613__B2 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6670_ _0174_ net52 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ _0844_ _0845_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ mod.registers.r7\[0\] _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4169__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3916__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _0717_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5483_ _2254_ _2373_ _2376_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5669__A2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4434_ _1402_ _1403_ _1313_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4365_ _1333_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6104_ _1999_ _2766_ _2806_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3316_ _3166_ _3168_ _3160_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1265_ _1070_ _0460_ _0452_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6035_ _2746_ mod.pc0\[7\] _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3451__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__B2 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A3 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6937_ _0035_ net175 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3604__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5378__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _0369_ net196 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5819_ _2598_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _0303_ net64 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3368__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3907__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3626__I _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__A2 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6844__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6994__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3536__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4323__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__B1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4150_ _1111_ _1112_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_110_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ mod.pc_2\[2\] _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4087__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_260 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_271 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_282 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_293 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _1627_ _1645_ _1385_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3598__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6722_ _0226_ net39 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3934_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5339__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3865_ mod.registers.r15\[10\] _0765_ _0766_ mod.registers.r12\[10\] _0835_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6653_ _0157_ net159 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5604_ mod.registers.r6\[11\] _2460_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _0515_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6584_ _3139_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ mod.registers.r5\[7\] _2405_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3365__A3 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4562__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5466_ mod.registers.r4\[3\] _2362_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3890__B _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4417_ _0949_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5397_ _2268_ _2315_ _2320_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6867__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4348_ _0828_ _0861_ _1253_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4277__I _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4078__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4279_ _1094_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6018_ _2736_ _1959_ _1965_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A1 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3825__B2 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5578__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4250__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3761__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4069__B2 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3816__B2 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A3 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__B2 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5746__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3694__C _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3650_ _0595_ _0599_ _0613_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A1 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3581_ _0530_ _0528_ _0539_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5320_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ mod.registers.r3\[11\] _0694_ _0879_ mod.registers.r7\[11\] _1172_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3504__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _1907_ _2136_ _1377_ _0984_ _2072_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_68_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4133_ _1047_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ mod.registers.r11\[6\] _3202_ _3194_ mod.registers.r10\[6\] mod.registers.r2\[6\]
+ _3190_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_84_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4480__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout42_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ _1388_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6705_ _0209_ net52 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3917_ _3172_ _3214_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4897_ mod.ldr_hzd\[15\] _1852_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3991__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6636_ _0140_ net142 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3848_ mod.registers.r4\[11\] _0419_ _3264_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4535__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _3118_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3779_ _0747_ _0433_ _0661_ _0563_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_164_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5518_ _2400_ _2389_ _2401_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6498_ _3087_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _2290_ _2349_ _2353_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4299__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3904__I _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout110 net125 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout132 net133 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout154 net156 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout165 net166 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout176 net179 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout187 net189 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout198 net199 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5799__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__I0 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4223__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4223__B2 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5566__I _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4403__C _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6598__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4526__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3734__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5250__B _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout177_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6203__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5962__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4765__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ _1228_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4380__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ mod.registers.r6\[1\] _0503_ _0515_ mod.registers.r12\[1\] _0672_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4682_ _1444_ _1456_ _1151_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3633_ _3198_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6421_ _1813_ _3033_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5714__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3725__B1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3564_ _3282_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6352_ _2985_ _2991_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5303_ _2178_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6283_ mod.des.des_dout\[18\] _2900_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3724__I _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3495_ _3173_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _2181_ _1910_ _2174_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _2107_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ mod.registers.r15\[5\] _0485_ _3208_ mod.registers.r14\[5\] _1086_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5096_ mod.pc_2\[8\] _2042_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6905__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4047_ _0482_ _0483_ mod.registers.r1\[7\] _1014_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4205__A1 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ mod.valid1 _2709_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4205__B2 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5953__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ mod.pc_2\[1\] _1046_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5705__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6619_ _0123_ net135 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4508__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5335__B _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__I _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6433__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4444__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4747__A2 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3707__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3544__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6928__CLK net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6970_ _0068_ net59 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _2421_ _2667_ _2670_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4986__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6188__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5852_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4199__B1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4803_ _1769_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5935__A1 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _2546_ _2579_ _2583_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4734_ _1437_ _1703_ _1243_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _1406_ _1362_ _1533_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_135_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _0687_ _2956_ _3024_ _2855_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3616_ mod.registers.r15\[5\] _0434_ _0436_ mod.registers.r12\[5\] _0586_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5163__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4596_ _1541_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6335_ _0636_ _2975_ _2979_ mod.instr\[12\] _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3547_ _0439_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4910__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6112__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ mod.instr\[14\] _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3478_ _0444_ _0445_ _0410_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5217_ _1786_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6197_ mod.pc_1\[10\] _2877_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4674__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5148_ _1907_ _2090_ _2105_ _3156_ _2106_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6415__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5079_ _1896_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6351__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__B2 mod.instr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3704__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__B1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3468__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4665__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6406__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5754__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3943__A3 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4450_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3401_ _3252_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4381_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6120_ _1925_ _2048_ _2051_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3332_ _3181_ _3167_ _3183_ _3184_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_98_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2722_ _2114_ _2117_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5002_ _1385_ _1621_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4959__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6953_ _0051_ net147 mod.ldr_hzd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ mod.registers.r13\[3\] _2656_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6884_ _0385_ net163 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ mod.registers.r11\[10\] _2613_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5908__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _2570_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5384__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4989__B _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _0497_ _0827_ _0841_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4592__B1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5664__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ _2431_ _2521_ _2523_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6333__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ _1095_ _1370_ _1548_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6333__B2 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4579_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__A1 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ mod.instr_2\[6\] _2968_ _2963_ mod.instr\[6\] _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6249_ _2918_ _2913_ _2919_ _2917_ _2911_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3912__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5839__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5072__B2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3622__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3359__I mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6773__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5574__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3689__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3310__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__I _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _3248_ _0916_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3613__A2 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3881_ _0777_ _0847_ _0849_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_149_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5620_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4023__C1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4169__A3 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5551_ _2267_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4502_ _1467_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5482_ mod.registers.r4\[9\] _2374_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _0525_ _0461_ _0592_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4341__A3 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4364_ _1205_ _0799_ _3262_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6103_ _2767_ _2805_ _2778_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3315_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _0578_ _0494_ _1069_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_99_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6034_ _2736_ _2032_ _2035_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout72_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6646__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__I _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _0034_ net162 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4801__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6867_ _0368_ net196 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5818_ _2538_ _2599_ _2605_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6798_ _0302_ net59 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3368__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3368__B2 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5749_ _2275_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5293__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6545__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4020__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4859__B2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3531__B2 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ _1033_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4087__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_250 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_261 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3834__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_272 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_283 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_294 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5479__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5036__B2 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__C1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0699_ _0710_ _3223_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3598__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6721_ _0225_ net50 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3598__B2 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3933_ _3230_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5339__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6652_ _0156_ net134 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6536__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ mod.registers.r9\[10\] _0751_ _0752_ mod.registers.r3\[10\] _0834_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _2425_ _2459_ _2463_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6583_ net17 mod.des.des_dout\[27\] _3137_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _0514_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3727__I _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5534_ _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3770__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5465_ _2194_ _2360_ _2365_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4416_ _0943_ _1380_ _1381_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_160_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5396_ mod.registers.r2\[11\] _2316_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4347_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _1033_ _1049_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4078__A2 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2728_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3825__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5027__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _0017_ net187 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3589__B2 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4250__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6527__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3761__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3761__B2 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5852__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6550__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3372__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A2 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5266__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6961__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4931__I _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3547__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout122_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _0540_ _0543_ _0546_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5250_ mod.des.des_dout\[24\] _2167_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3504__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4201_ _1168_ _1169_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3504__B2 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__B1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5181_ _1907_ _2136_ _1435_ _1001_ _2072_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_96_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4132_ _1050_ _1073_ _1096_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__A1 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4480__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _1932_ _1604_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6704_ _0208_ net92 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ _0880_ _0881_ _0883_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4896_ _1848_ _1860_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6635_ _0139_ net141 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3991__B2 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3847_ mod.registers.r11\[11\] _0505_ _0412_ mod.registers.r2\[11\] _0817_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6834__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6566_ _3128_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ mod.registers.r15\[12\] _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4535__A3 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5517_ mod.registers.r5\[3\] _2391_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ mod.des.des_dout\[9\] net7 _3085_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5448_ mod.registers.r3\[14\] _2350_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5496__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout100 net110 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout111 net115 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5379_ _2303_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout122 net123 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout133 net144 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout144 net145 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout155 net156 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout166 net167 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout177 net179 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout188 net189 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__I1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6008__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__I _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5971__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3982__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3734__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3734__B2 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4926__I _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6707__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4214__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _1247_ _1706_ _1707_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3701_ mod.registers.r13\[1\] _0520_ _3272_ mod.registers.r8\[1\] _0671_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4681_ _1279_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6420_ _3034_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3632_ _3194_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3725__A1 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3725__B2 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ mod.funct7\[0\] _2989_ _2986_ mod.instr\[18\] _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3563_ mod.registers.r8\[7\] _0531_ _0532_ mod.registers.r10\[7\] _0533_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6282_ mod.instr\[18\] _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3494_ _3265_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5233_ mod.pc_2\[1\] _2182_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5164_ _1727_ _1737_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ mod.registers.r8\[5\] _3204_ _3198_ mod.registers.r9\[5\] _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _1970_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ mod.registers.r3\[7\] _1013_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4453__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _2712_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4205__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5402__A1 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4948_ _1206_ _3259_ _1077_ _3263_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4504__C _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4879_ _0490_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6618_ _0122_ net138 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5181__A3 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4141__A1 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__I _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6433__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4444__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6197__A2 _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3707__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3707__B2 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6201__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A2 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4683__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3560__I mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5632__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ mod.registers.r13\[9\] _2668_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6188__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4199__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _1182_ _1397_ _1641_ _1330_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4199__B2 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5782_ mod.registers.r10\[6\] _2580_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5935__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ _1442_ _1682_ _1675_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5148__B1 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _1541_ _1612_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_135_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5699__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ mod.ri_3 _2867_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3615_ _0581_ _0582_ _0583_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_128_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6360__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3735__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ _1357_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6334_ _2978_ _2980_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3546_ mod.registers.r15\[6\] _0514_ _0515_ mod.registers.r12\[6\] _0516_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4910__A3 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _2930_ _2925_ _2931_ _2929_ _2923_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6112__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5950__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4123__A1 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6196_ _2872_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5871__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4674__A2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5171__B _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3470__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5147_ _1171_ _1176_ _1929_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _1909_ _1511_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input15_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4029_ mod.registers.r3\[14\] _0959_ _0960_ mod.registers.r2\[14\] _0999_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3634__B1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6351__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4114__A1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5862__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3380__I _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__B _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3555__I _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout202_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4353__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4380_ _0621_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ mod.instr_2\[14\] _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _2759_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5001_ _1949_ _1967_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__B1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5605__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _0050_ net152 mod.ldr_hzd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3616__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _2396_ _2654_ _2659_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6883_ _0384_ net155 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _2554_ _2612_ _2615_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5908__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5765_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4716_ _1317_ _1409_ _1592_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5696_ mod.registers.r8\[12\] _2522_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4647_ _1074_ _1337_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3465__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4578_ _0930_ _0932_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6317_ _2961_ _2969_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3529_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ mod.des.des_dout\[9\] _2909_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6179_ _2860_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3855__B1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6021__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6918__CLK net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4583__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5076__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3375__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A2 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6088__A1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3846__B1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout152_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3880_ _0846_ _0632_ mod.registers.r8\[8\] _0638_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A1 _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4023__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__C2 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5550_ _2425_ _2418_ _2426_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4501_ _0925_ _1410_ _1414_ _1469_ _1470_ _1315_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_157_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _2245_ _2373_ _2375_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4432_ _1401_ _1310_ _0576_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4363_ _0692_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6079__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6102_ _2801_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3314_ mod.instr_2\[16\] _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_112_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _0625_ _0680_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4629__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _2743_ _2748_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5005__I mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0033_ net175 mod.ri_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6866_ _0367_ net196 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ mod.registers.r11\[3\] _2601_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _0301_ net64 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5675__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3368__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _2558_ _2551_ _2559_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5679_ _2408_ _2509_ _2512_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__A1 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5817__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3828__B1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6740__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4308__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3531__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4087__A3 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_240 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6365__B _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_251 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_262 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3834__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_273 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_284 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6084__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_295 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6233__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4981_ _1931_ _1948_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4244__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__C2 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _0224_ net92 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3598__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3932_ _0457_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6651_ _0155_ net138 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3863_ _0829_ _0830_ _0831_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6536__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ mod.registers.r6\[10\] _2460_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6582_ _3138_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3794_ _0760_ _0761_ _0762_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_118_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5533_ _2235_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3770__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5464_ mod.registers.r4\[2\] _2362_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4415_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5395_ _2261_ _2315_ _2319_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6613__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4346_ _0801_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4277_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6016_ _2733_ _2735_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6472__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6918_ _0016_ net154 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _0350_ net192 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3761__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4171__C1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6463__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4484__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4433__B _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6636__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout115_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ mod.registers.r6\[11\] _0700_ _0889_ mod.registers.r13\[11\] _1170_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3504__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _2107_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6786__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _1097_ _1049_ _1098_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_122_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _1030_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _1385_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6703_ _0207_ net55 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ mod.registers.r15\[4\] _0884_ _0600_ mod.registers.r6\[4\] _0603_ mod.registers.r9\[4\]
+ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_4895_ _1861_ _1863_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3846_ mod.registers.r14\[11\] _0502_ _0503_ mod.registers.r6\[11\] _0816_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3991__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6634_ _0138_ net140 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6565_ mod.des.des_dout\[20\] net5 _3124_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3777_ mod.registers.r12\[12\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5516_ _2399_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3743__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6496_ _3086_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5447_ _2284_ _2349_ _2352_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5496__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout101 net104 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5378_ _2301_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout134 net137 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4329_ _0991_ _1296_ _1297_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xfanout145 net146 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout156 net157 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout167 net168 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout178 net179 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout189 net194 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4518__B _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__I2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3982__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5863__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3734__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4998__B2 _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4942__I _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3558__I _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ mod.registers.r1\[1\] _0521_ _0412_ mod.registers.r2\[1\] _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _1648_ _1649_ _1128_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5175__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3631_ mod.registers.r6\[2\] _0600_ _3189_ mod.registers.r5\[2\] mod.registers.r2\[2\]
+ _3191_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6350_ _2985_ _2990_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3562_ _3278_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3725__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5301_ mod.des.des_dout\[29\] _2188_ _2240_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_127_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ _2942_ _2937_ _2943_ _2941_ _2935_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3493_ _0454_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5232_ _1793_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3489__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _1196_ _1199_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6427__A1 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ mod.registers.r4\[5\] _0465_ _3194_ mod.registers.r10\[5\] _1084_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ _1909_ _1674_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4338__B _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4045_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6801__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _1789_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4878_ mod.instr_2\[6\] _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6617_ _0121_ net135 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6951__CLK net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ _0791_ _0796_ _0797_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_146_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3716__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ mod.des.des_counter\[2\] _1906_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6479_ mod.des.des_dout\[1\] net17 _3075_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4141__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3707__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__I _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4132__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6824__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__B1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5850_ _2357_ _2624_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _1180_ _1670_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4199__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A1 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _2544_ _2579_ _2582_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4732_ _1256_ _1678_ _1700_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ _0989_ _1538_ _1345_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5148__B2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4621__B _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _3021_ _3022_ _3023_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5699__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3614_ mod.registers.r4\[5\] _0418_ _3236_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4594_ _0989_ _1316_ _1341_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3545_ _0436_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6333_ _1808_ _2975_ _2979_ mod.instr\[11\] _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4910__A4 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6264_ mod.des.des_dout\[13\] _2921_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout95_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3476_ _0444_ _0445_ _3281_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4123__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _2066_ _2876_ _2879_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5146_ _2101_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5871__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3882__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _2037_ _2038_ _2039_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5623__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4028_ mod.registers.r15\[14\] _0964_ _0968_ mod.registers.r8\[14\] _0998_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3634__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3634__B2 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4434__I0 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5979_ net11 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6503__S _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4898__C2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3570__B1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6847__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6997__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3928__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4050__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6212__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4889__B1 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5550__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4353__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3571__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _3225_ _1950_ _1966_ _1904_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__B2 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5605__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7002__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _0049_ net150 mod.ldr_hzd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5498__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3616__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3616__B2 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ mod.registers.r13\[2\] _2656_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6882_ _0383_ net151 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5833_ mod.registers.r11\[9\] _2613_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4041__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6318__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4715_ _1436_ _1680_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3746__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5695_ _2503_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4646_ _1518_ _1269_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _1076_ _1099_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3552__B1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _2967_ _2968_ _2963_ mod.instr\[5\] _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_131_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ _0457_ _3257_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3459_ _3289_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6247_ mod.instr\[9\] _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3855__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3855__B2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _3225_ _2074_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__A1 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5780__A1 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5532__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3543__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6188__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5092__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3605__B _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A3 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3846__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3846__B2 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5599__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6260__A2 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__I mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout145_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4023__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _1403_ _1413_ _0496_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5480_ mod.registers.r4\[8\] _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4431_ _0667_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5523__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__B1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4362_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6101_ _1998_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3313_ _3161_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4397__I _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4293_ _1260_ _1261_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _2746_ mod.pc0\[6\] _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3837__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout58_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6117__I _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _0032_ net175 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4262__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _0366_ net197 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5816_ _2536_ _2599_ _2604_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6796_ _0300_ net120 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5747_ mod.registers.r9\[11\] _2552_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4565__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ mod.registers.r8\[5\] _2510_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5514__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0576_ _0592_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3828__B2 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4253__A1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6471__B _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3386__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3764__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5505__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4010__I _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4945__I _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_230 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4492__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_241 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_252 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_263 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_274 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_285 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_296 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6233__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _3225_ _1933_ _1947_ _1904_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4244__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4244__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3931_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5776__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _0154_ net138 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ mod.registers.r4\[10\] _0420_ _3265_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5601_ _2422_ _2459_ _2462_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5744__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ net16 mod.des.des_dout\[26\] _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3793_ mod.registers.r4\[13\] _0738_ _3238_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5532_ _2411_ _2404_ _2412_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ _2186_ _2360_ _2364_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3770__A3 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__S _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4414_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5394_ mod.registers.r2\[10\] _2316_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0809_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4276_ _0940_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6908__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2734_ mod.pc0\[2\] _2731_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4855__I mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6917_ _0015_ net156 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4786__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6848_ _0349_ net198 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _0283_ net136 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3934__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4171__B1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__C2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6463__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3737__B1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4005__I _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3844__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__A1 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4701__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ _1076_ _1099_ _1075_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4061_ _1029_ _1022_ _1026_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4217__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _0599_ _0613_ _3223_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _0206_ net49 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3914_ _0485_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4894_ mod.ldr_hzd\[6\] _1858_ _1854_ mod.ldr_hzd\[5\] _1851_ mod.ldr_hzd\[7\] _1864_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5717__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6633_ _0137_ net140 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3845_ mod.registers.r8\[11\] _0531_ _0500_ mod.registers.r10\[11\] _0815_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3728__B1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _3127_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3776_ _0521_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5515_ _2198_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6495_ mod.des.des_dout\[8\] net6 _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3754__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5446_ mod.registers.r3\[13\] _2350_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5377_ _2199_ _2302_ _2308_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout102 net104 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3900__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout135 net137 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4328_ _1296_ _1297_ _0992_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout146 net204 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout157 net158 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3703__B _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout168 net169 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout179 net183 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4259_ _1226_ _1201_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4456__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6880__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__B2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__I3 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4208__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6381__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6040__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__S _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3742__I0 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4444__B _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3839__I _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3630_ _3185_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5175__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6372__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3561_ _3271_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3574__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _2213_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6124__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6280_ mod.des.des_dout\[17\] _2933_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _0461_ _0453_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _1793_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4686__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3489__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _2109_ _2119_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4150__A3 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__B _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4113_ mod.registers.r12\[5\] _0887_ _3185_ mod.registers.r6\[5\] _1083_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5093_ _1908_ _2040_ _2053_ _0001_ _2054_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _3166_ _3216_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout40_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6125__I _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4946_ _1789_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4877_ _1838_ _1841_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_138_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _0120_ net130 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ mod.registers.r8\[15\] _0729_ _0765_ mod.registers.r15\[15\] _0798_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6363__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ _2441_ _3112_ _3117_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3759_ _3272_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4913__A2 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6478_ _3076_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _2229_ _2337_ _2341_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4677__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__B _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__I _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6776__CLK net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6354__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6354__B2 mod.instr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3394__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__B2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__B _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__B1 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout175_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _1181_ _1484_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ mod.registers.r10\[5\] _2580_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4731_ _1700_ _1256_ _1678_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _0925_ _1561_ _1630_ _1306_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__5148__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _2715_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3613_ mod.registers.r11\[5\] _3291_ _0411_ mod.registers.r2\[5\] _0583_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4593_ _1559_ _1562_ _1327_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6332_ _2950_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3544_ _0434_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ mod.instr\[13\] _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3475_ _0426_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ _2142_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6194_ mod.pc_1\[9\] _2877_ _2873_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout88_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4349__B _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ mod.pc0\[11\] _1892_ _1901_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3882__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _1008_ _1020_ _1985_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5959__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4027_ mod.registers.r6\[14\] _0966_ _0967_ mod.registers.r5\[14\] _0997_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3634__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4831__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6799__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3479__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _2441_ _2700_ _2705_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4434__I1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _1884_ _1889_ _1895_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5694__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5139__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3570__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3570__B2 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3942__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6474__B _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3389__I _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4035__C1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A3 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__B _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5066__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__CLK net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6950_ _0048_ net149 mod.ldr_hzd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3616__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ _2393_ _2654_ _2658_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6881_ _0382_ net151 mod.instr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _2550_ _2612_ _2614_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5763_ _2299_ _2499_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4632__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4041__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4714_ _1243_ _1683_ _1433_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6318__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _2501_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4645_ _1518_ _1514_ _1241_ _0940_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5019__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3927__I0 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _1306_ _1544_ _1545_ _1309_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3552__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _2955_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3552__B2 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3527_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3762__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6246_ _2915_ _2913_ _2916_ _2917_ _2911_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3458_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6177_ _2857_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3389_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3855__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _2084_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5057__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _1037_ _1042_ _1985_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4804__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4280__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6313__I _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6309__A1 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__B2 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5780__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3791__B2 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5532__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3543__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4768__I _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3543__B2 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__I0 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6964__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5048__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4008__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4452__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6223__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout138_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _0726_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__B _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__B2 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__I _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _0917_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3582__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6100_ _2802_ _2769_ mod.pc\[5\] _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3312_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4292_ _0723_ _0666_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _2736_ _2016_ _2019_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__I _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6933_ _0031_ net164 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4262__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _0365_ net195 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5815_ mod.registers.r11\[2\] _2601_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6795_ _0299_ net117 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3757__I mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _2267_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ _2403_ _2509_ _2511_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4628_ _1313_ _0555_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__CLK net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3525__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4559_ _1320_ _1354_ _1344_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__A4 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ _2891_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3828__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5212__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4253__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5753__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3764__B2 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6199__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3516__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_231 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_242 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6218__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_253 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_264 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_275 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_286 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_297 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3930_ _0878_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5278__B _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ mod.registers.r11\[10\] _3292_ _0413_ mod.registers.r2\[10\] _0831_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3577__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5600_ mod.registers.r6\[9\] _2460_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6580_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5744__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3792_ mod.registers.r11\[13\] _0735_ _0736_ mod.registers.r2\[13\] _0762_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ mod.registers.r5\[6\] _2405_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ mod.registers.r4\[1\] _2362_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3507__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4413_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5393_ _2254_ _2315_ _2318_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4180__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ _1309_ _1312_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _1240_ _1243_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ _2728_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout70_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _0014_ net149 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6847_ _0348_ net190 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _0282_ net136 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5729_ _2228_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4171__B2 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4474__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3521__I1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3682__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3737__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__B2 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4956__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ _1022_ _1026_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4870__C1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__A1 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _1908_ _1910_ _1928_ _0001_ _1930_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__5965__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6701_ _0205_ net54 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3913_ mod.registers.r5\[4\] _0882_ _0706_ mod.registers.r8\[4\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3976__A1 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ mod.ldr_hzd\[4\] _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6632_ _0136_ net126 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3844_ _0557_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3728__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ mod.des.des_dout\[19\] net4 _3124_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3728__B2 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3775_ _0520_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4640__B _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6390__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5514_ _2397_ _2389_ _2398_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ _3074_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5445_ _2276_ _2349_ _2351_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4153__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ mod.registers.r2\[3\] _2304_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout103 net104 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3900__A1 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout114 net115 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4327_ _1003_ _1232_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout125 net145 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3900__B2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout136 net139 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout147 net150 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout158 net169 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _1221_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout169 net185 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5653__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ mod.registers.r14\[10\] _0891_ _0703_ mod.registers.r9\[10\] mod.registers.r2\[10\]
+ _0893_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4534__C _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4106__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3719__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6908__D _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3742__I1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4447__A2 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A2 _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout120_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout218_I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ mod.pc_2\[7\] _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_142_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3491_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5230_ _2164_ _2177_ _2180_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4135__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5291__B _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _1985_ _1218_ _2118_ _1969_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ _1079_ _1080_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ _1131_ _1142_ _1929_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5635__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _3209_ _3217_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ mod.valid0 _2709_ _2151_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3949__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4945_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4071__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _1842_ _1843_ _1844_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3827_ mod.registers.r11\[15\] _0735_ _0738_ mod.registers.r4\[15\] _0736_ mod.registers.r2\[15\]
+ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6615_ _0119_ net131 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3765__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6546_ mod.registers.r15\[15\] _3113_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3758_ _3266_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6477_ mod.des.des_dout\[0\] net16 _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5980__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3689_ mod.registers.r9\[3\] _0544_ _0545_ mod.registers.r3\[3\] _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4126__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ mod.registers.r3\[6\] _2338_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ mod.des.des_dout\[36\] _2220_ _2292_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__3885__B1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4365__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__S _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5865__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3624__B _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3628__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5093__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__B2 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__B _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout168_I net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _1437_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__B1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _1318_ _1321_ _0626_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6400_ _1886_ _1798_ _3249_ _2858_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3612_ mod.registers.r14\[5\] _3282_ _3286_ mod.registers.r6\[5\] _0582_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _0692_ _1560_ _1561_ _0626_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _2759_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3543_ mod.registers.r9\[6\] _0511_ _0512_ mod.registers.r3\[6\] _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6262_ _2927_ _2925_ _2928_ _2929_ _2923_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3474_ _0425_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5856__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6193_ _2050_ _2876_ _2878_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3867__B1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5144_ _2102_ _2041_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _1987_ _2024_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3619__B1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5084__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _0993_ _0994_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__A2 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5040__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6033__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ mod.registers.r14\[15\] _2701_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _1893_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _0640_ _1816_ _1821_ _0848_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4898__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _3094_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3570__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5075__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__B1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__C2 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__CLK net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4050__A3 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4889__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__I mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A4 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5066__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5900_ mod.registers.r13\[1\] _2656_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _0381_ net151 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6015__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5831_ mod.registers.r11\[8\] _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ _2568_ _2561_ _2569_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4041__A3 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4713_ _1442_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _2428_ _2515_ _2520_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6318__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _1609_ _1610_ _1612_ _1566_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_135_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3927__I1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4575_ _1468_ _1501_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3552__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3526_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6314_ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _2891_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3457_ _0424_ _3269_ _0425_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ _1962_ _2859_ _2866_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3388_ _3227_ _3229_ _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5127_ mod.pc0\[10\] _1922_ _1923_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6254__B2 _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ _1987_ _2007_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4009_ mod.registers.r14\[15\] _0977_ _0978_ mod.registers.r7\[15\] _0979_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__A3 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3791__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3953__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3543__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__I1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5296__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5048__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4733__B _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5220__A2 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6639__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout200_I net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1328_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3311_ _3160_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4291_ _0807_ _0650_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ _2722_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _0030_ net165 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6863_ _0364_ net188 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ _2534_ _2599_ _2603_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6794_ _0298_ net117 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5211__A2 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5745_ _2556_ _2551_ _2557_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4970__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ mod.registers.r8\[4\] _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4627_ _0593_ _0860_ _0875_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3773__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__C1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _1318_ _1321_ _1406_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3509_ mod.registers.r12\[1\] _0476_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4489_ _1228_ _1222_ _1458_ _1285_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6228_ mod.des.des_dout\[4\] _2896_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6159_ _2850_ _2852_ _2818_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3948__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3764__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3516__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6466__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_232 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_243 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_254 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_265 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_276 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_287 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4019__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_298 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3452__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3858__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout150_I net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3860_ mod.registers.r14\[10\] _0732_ _0733_ mod.registers.r6\[10\] _0830_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ mod.registers.r14\[13\] _3283_ _3287_ mod.registers.r6\[13\] _0761_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5461_ _2177_ _2360_ _2363_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4412_ _0942_ _0932_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5392_ mod.registers.r2\[9\] _2316_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ _0923_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4180__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__B2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _1239_ _1004_ _1238_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_140_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _2726_ _1947_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout63_I net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _0013_ net81 mod.instr_2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3768__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _0347_ net178 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5983__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _0281_ net134 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3989_ _3165_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5728_ _2544_ _2541_ _2545_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5659_ _2149_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4171__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3682__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3682__B2 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6229__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6827__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4870__C2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__B _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _0470_ _0488_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6700_ _0204_ net113 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3912_ _3188_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3976__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4892_ _1856_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5178__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _0135_ net130 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3843_ _0556_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3728__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6562_ _3126_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3774_ mod.registers.r7\[12\] _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5513_ mod.registers.r5\[2\] _2391_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6493_ _3084_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5444_ mod.registers.r3\[12\] _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4153__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5350__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _2194_ _2302_ _2307_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout104 net109 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout115 net124 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3900__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4326_ _1287_ _1295_ _1236_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_59_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout126 net133 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_141_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout137 net139 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout148 net150 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout159 net160 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4257_ _1226_ _1201_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5653__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4188_ mod.registers.r6\[10\] _0700_ _0705_ mod.registers.r11\[10\] _1158_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3664__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3498__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6829_ _0000_ _0004_ net218 mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4144__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3352__B1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5892__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3407__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4907__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5580__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3490_ _0455_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4135__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _2114_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__B2 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ mod.registers.r5\[5\] _3188_ _3211_ mod.registers.r13\[5\] _1081_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5091_ _2049_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5635__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4042_ _0951_ _3216_ mod.registers.r4\[7\] _1010_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5993_ _2710_ _2714_ _2716_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1911_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4071__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4071__B2 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4875_ _1802_ _1834_ _1835_ _1810_ _1836_ _1804_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_32_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6422__I _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6614_ _0118_ net130 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3826_ _0792_ _0793_ _0794_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6545_ _2438_ _3112_ _3116_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5571__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ mod.pc_2\[12\] _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ _3074_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3688_ mod.registers.r7\[3\] _0548_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5427_ _2218_ _2337_ _2340_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5323__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3781__I _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5358_ _2226_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3885__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3885__B2 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ _0873_ _1124_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5289_ _1935_ _2208_ _2226_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5501__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4062__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3956__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6332__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4365__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6672__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3573__B1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4117__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3691__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5865__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4736__B _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3628__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3628__B2 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6507__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5411__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__B2 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4660_ _1628_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3611_ mod.registers.r8\[5\] _3271_ _3278_ mod.registers.r10\[5\] _0581_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5553__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _0666_ _1251_ _0667_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _2971_ _2977_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3542_ _0430_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6398__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4108__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ net13 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3473_ mod.registers.r5\[0\] _0440_ _0442_ mod.registers.r7\[0\] _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5212_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6192_ mod.pc_1\[8\] _2877_ _2873_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3867__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3867__B2 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5143_ mod.pc\[11\] _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ _1969_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3619__B2 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ mod.registers.r11\[14\] _0974_ _0980_ mod.registers.r13\[14\] _0995_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4292__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _2438_ _2700_ _2704_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4044__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5792__A1 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3776__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _1823_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3809_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6592__I0 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4789_ _1281_ _1650_ _1741_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _3092_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _1802_ _3058_ _3059_ _3044_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4035__B2 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__I0 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6011__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout180_I net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5830_ _2600_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ mod.registers.r9\[15\] _2562_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4577__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4041__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4712_ _1518_ _1096_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5692_ mod.registers.r8\[11\] _2516_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6574__I0 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _1501_ _1419_ _0776_ _0803_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3537__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ _1312_ _1319_ _0593_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1861_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3525_ _0464_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6244_ mod.des.des_dout\[8\] _2909_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ mod.instr_2\[10\] _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4501__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ mod.pc_1\[3\] _2861_ _2864_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3387_ _3233_ _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _2085_ _1897_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4376__B _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6254__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _1969_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4008_ _3170_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _2680_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A1 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6565__I0 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4740__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__B1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__I _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6860__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3767__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__I mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3310_ _3161_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4290_ _1062_ _1063_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4196__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6236__A2 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _0029_ net165 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4798__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _0363_ net196 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5813_ mod.registers.r11\[1\] _2601_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5747__A1 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _0297_ net118 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4215__I _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ mod.registers.r9\[10\] _2552_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _2503_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4970__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _1327_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6733__CLK net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4183__C2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ _1524_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4722__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3508_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4488_ _1444_ _1456_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6227_ mod.instr\[4\] _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3439_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4486__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6883__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6158_ _2850_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _1109_ _1120_ _1929_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ _2783_ _2785_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4238__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4410__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4961__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput30 net30 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_233 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_244 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_255 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_266 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_277 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_288 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5977__A1 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_299 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6606__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3452__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout143_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3790_ mod.registers.r8\[13\] _3273_ _3279_ mod.registers.r10\[13\] _0760_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6250__I mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ mod.registers.r4\[0\] _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0943_ _1377_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5901__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2245_ _2315_ _2317_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _0527_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4919__B mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4273_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4468__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6012_ _2730_ _1928_ _2732_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

