* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5968__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout56_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _0012_ net143 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4640__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6845_ _0346_ net153 mod.pc0\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6776_ _0280_ net67 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3988_ _0951_ _0954_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_22_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ mod.registers.r9\[5\] _2542_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6160__I _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _2442_ _2492_ _2497_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4609_ _0948_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5589_ _2403_ _2453_ _2455_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3903__B1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6448__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5504__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6629__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3682__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4564__B _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4698__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4739__B _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4870__B2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _3153_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3911_ mod.registers.r3\[4\] _3165_ _0697_ mod.registers.r1\[4\] _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4891_ mod.instr_2\[5\] _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6630_ _0134_ net87 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3842_ _0801_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5178__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6561_ mod.des.des_dout\[18\] net3 _3124_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3773_ _0518_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5512_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6492_ mod.des.des_dout\[7\] net5 _3080_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4138__B1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5443_ _2331_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5350__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ mod.registers.r2\[2\] _2304_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout105 net107 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout127 net128 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout138 net140 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4256_ _0773_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ mod.registers.r1\[10\] _0697_ _0980_ mod.registers.r13\[10\] _1157_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4861__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3664__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6921__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4613__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ _0332_ net44 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6759_ _0263_ net67 mod.registers.r10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__B _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__A3 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3352__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3352__B2 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__I0 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3407__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4907__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4135__A3 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5332__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ mod.registers.r3\[5\] _0471_ _0466_ mod.registers.r1\[5\] _3201_ mod.registers.r11\[5\]
+ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_110_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ mod.pc0\[8\] _1892_ _1901_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5096__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6944__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4041_ _3215_ _3168_ mod.registers.r8\[7\] _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5992_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _1787_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ _1807_ _1832_ _1113_ _0711_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6613_ _0117_ net89 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3825_ mod.registers.r9\[15\] _0751_ _0730_ mod.registers.r10\[15\] _0795_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ mod.registers.r15\[14\] _3113_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3756_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5571__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ mod.des.des_counter\[0\] mod.des.des_counter\[1\] mod.des.des_counter\[2\]
+ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3687_ mod.registers.r5\[3\] _0547_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5426_ mod.registers.r3\[5\] _2338_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6520__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5357_ _0958_ _2224_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3885__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0840_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5288_ mod.pc_2\[7\] _2221_ _2224_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4239_ mod.registers.r4\[12\] _0971_ _0972_ mod.registers.r10\[12\] _1209_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4561__C _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5011__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4133__I _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3573__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3573__B2 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__A2 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6967__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3628__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4053__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5250__A1 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3610_ mod.pc_2\[5\] _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4590_ _1308_ _1311_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5553__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _0427_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ mod.des.des_dout\[12\] _2921_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5305__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3472_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3316__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _2150_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6191_ _2857_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3867__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _1924_ _2091_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _2032_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4024_ mod.registers.r14\[14\] _0977_ _0978_ mod.registers.r7\[14\] _0981_ mod.registers.r9\[14\]
+ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4292__A2 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ mod.registers.r14\[14\] _2701_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _1824_ _1806_ _0661_ _1825_ _0429_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4788_ _1720_ _1727_ _1737_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__6592__I1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _2413_ _3100_ _3105_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3739_ mod.registers.r14\[3\] _0607_ _0608_ mod.registers.r13\[3\] _0708_ _0709_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _2716_ _3062_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5409_ _2150_ _2327_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6389_ _2075_ _3009_ _3015_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__I _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5480__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4035__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3546__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__B2 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A1 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3849__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__B _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6518__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4274__A2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout173_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__B1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6253__I _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ _2295_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3785__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _1098_ _1100_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3785__B2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _2425_ _2515_ _2519_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4642_ _0900_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4329__A3 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6574__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3537__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3537__B2 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4573_ _1531_ _1536_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6312_ _2961_ _2965_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3524_ _3254_ _0470_ _0488_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6243_ mod.instr\[8\] _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3455_ mod.instr_2\[11\] _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout86_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6174_ _1944_ _2859_ _2865_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3386_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ mod.pc\[10\] _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6428__I _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _2016_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5462__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ _0607_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3473__B1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3787__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6163__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _2413_ _2688_ _2693_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _1826_ _1822_ _1824_ _1825_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5889_ mod.registers.r12\[14\] _2647_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3528__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__B2 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__C _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__I0 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5756__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6022__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6181__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__A3 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6685__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6930_ _0028_ net183 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _0362_ net186 mod.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ _2527_ _2599_ _2602_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6792_ _0296_ net67 mod.registers.r12\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3400__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5747__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5743_ _2260_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _2501_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _1350_ _1591_ _1593_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_129_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4183__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _0593_ _1353_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4183__B2 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3930__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ _3181_ _3162_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _1128_ _1151_ _1274_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_89_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _2899_ _2901_ _2902_ _2892_ _2898_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3438_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5683__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _2851_ _2132_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5062__I _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3369_ _3192_ _3200_ _3205_ _3221_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _2041_ _2065_ _2068_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6088_ _1959_ _2790_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5435__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4238__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _1989_ _2003_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6107__B mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5738__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4410__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput20 net20 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4477__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_223 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_234 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_245 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_256 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5426__A1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_267 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_278 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_289 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3988__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4316__I _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout136_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4410_ _0992_ _1377_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5390_ mod.registers.r2\[8\] _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4341_ _0757_ _0861_ _0650_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__C _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4468__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _2723_ mod.pc0\[1\] _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3676__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__C1 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5968__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__A1 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _0011_ net142 mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _0345_ net154 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ _0279_ net66 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3987_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6393__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5726_ _2217_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3600__B1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5657_ mod.registers.r7\[15\] _2493_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4156__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6850__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ _3250_ _1558_ _1571_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5588_ mod.registers.r6\[4\] _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3903__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ _0918_ _1505_ _1508_ _1149_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5656__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3305__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4631__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4136__I _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6552__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__B _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4395__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4147__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4698__A2 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5647__A1 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__A3 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4474__C _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6072__A1 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6723__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3425__A3 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3910_ mod.registers.r7\[4\] _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _1855_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3841_ _0622_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6261__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _3125_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3772_ mod.registers.r5\[12\] _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5511_ _2193_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6491_ _3083_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4138__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _2329_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4138__B2 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ _2186_ _2302_ _2306_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _1288_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout106 net107 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout117 net118 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5638__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout128 net151 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout139 net140 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4255_ _1184_ _1190_ _1204_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4310__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ _1153_ _1154_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A2 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3821__B1 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6827_ _0331_ net44 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3795__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6758_ _0262_ net71 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6689_ _0193_ net99 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__B _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5515__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__A4 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3352__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__I1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__B1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5801__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4604__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6896__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4907__A3 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A1 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5096__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4040_ _0476_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6256__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2706_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1389_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6205__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4873_ _1826_ _1834_ _1835_ _1822_ _1825_ _1832_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_6612_ _0116_ net146 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3824_ mod.registers.r1\[15\] _0746_ _0431_ mod.registers.r3\[15\] _0794_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3406__I0 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5020__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6543_ _2435_ _3112_ _3115_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3755_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6619__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _3072_ _3073_ _2789_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3686_ _0652_ _0653_ _0654_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2205_ _2337_ _2339_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5356_ _2168_ _2107_ _1377_ _2273_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_114_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _1161_ _1164_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5287_ _2181_ _2024_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__A2 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _1136_ _1206_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ mod.registers.r3\[8\] _1013_ _1015_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4598__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5245__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5078__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__B1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5250__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3368__C _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout216_I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ _0501_ _0504_ _0507_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6911__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3471_ _0415_ _0416_ _3289_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5210_ _2155_ _2157_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6190_ _2867_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__I _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5141_ _2092_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5072_ mod.pc0\[7\] _1960_ _1961_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ mod.registers.r4\[14\] _0971_ _0975_ mod.registers.r1\[14\] _0972_ mod.registers.r10\[14\]
+ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_38_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6861__D _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5974_ _2435_ _2700_ _2703_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4662__C _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__A2 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4856_ mod.ldr_hzd\[7\] _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3807_ _0498_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4787_ _1743_ _1747_ _1748_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ mod.registers.r15\[7\] _3101_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4752__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3738_ _0660_ _3213_ _3214_ _3218_ _0662_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ _1810_ _3058_ _3059_ _3041_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3669_ _0424_ _0636_ mod.registers.r4\[2\] _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3307__A2 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _2160_ _2298_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6388_ mod.pc_1\[10\] _3010_ _3012_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ mod.registers.r1\[12\] _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _0107_ net205 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__B _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3794__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6934__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3546__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6248__A1 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3482__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__B2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ _1678_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3785__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4982__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5690_ mod.registers.r8\[10\] _2516_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4641_ _0878_ _1341_ _0716_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3537__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4572_ _0900_ _1537_ _1540_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6311_ mod.instr_2\[4\] _2958_ _2963_ mod.instr\[4\] _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3523_ _0489_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6242_ _2912_ _2913_ _2914_ _2905_ _2911_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3454_ _3267_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3385_ _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6173_ mod.pc_1\[2\] _2861_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4657__C _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _1914_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ mod.pc0\[6\] _1960_ _1961_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4006_ mod.registers.r11\[15\] _0974_ _0975_ mod.registers.r1\[15\] _0976_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5462__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3473__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3473__B2 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6957__CLK net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ mod.registers.r14\[7\] _2689_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1820_ _1819_ _1818_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_21_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5888_ _2564_ _2646_ _2649_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4839_ _1808_ _0445_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4725__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3528__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3308__I mod.instr_2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4489__B1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5150__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3700__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__C1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3464__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3767__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4602__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4716__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__C1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6529__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5444__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6492__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _0361_ net189 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5811_ mod.registers.r11\[0\] _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4404__B1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _0295_ net66 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5742_ _2554_ _2551_ _2555_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5673_ _2400_ _2502_ _2508_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4624_ _0691_ _0808_ _0790_ _0800_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3915__C1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4183__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _0529_ _0681_ _0839_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3506_ _3175_ _3217_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3930__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4486_ _1448_ _1453_ _1454_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6225_ mod.des.des_dout\[3\] _2896_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3437_ _3267_ _3269_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6156_ _2130_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3368_ mod.registers.r14\[0\] _3208_ _3211_ mod.registers.r13\[0\] _3220_ _3221_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_97_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3694__B2 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5107_ _2066_ _1891_ _2067_ _2041_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6087_ _2782_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3299_ _0000_ mod.des.des_counter\[1\] _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6483__I1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5038_ _3223_ _1990_ _2002_ _1904_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _0087_ net211 mod.des.des_dout\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3749__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4174__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3685__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_224 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_235 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_246 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_257 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_268 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_279 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout129_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ _1059_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6259__I mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4271_ _0908_ _0910_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6311__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ _2140_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4873__B1 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4873__C2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3428__A1 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6912_ _0010_ net143 mod.instr_2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3979__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3411__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A3 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6843_ _0344_ net155 mod.pc0\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4928__A1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ _0278_ net72 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3986_ _0955_ _0952_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _2540_ _2541_ _2543_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3600__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5338__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3600__B2 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5656_ _2439_ _2492_ _2496_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4156__A2 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _1572_ _1556_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5587_ _2447_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4538_ _1506_ _0934_ _1507_ _1484_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3903__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__B1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4469_ _1337_ _1251_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5656__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _2717_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _2828_ _2827_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6118__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4919__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4395__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A1 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A2 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A3 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3425__A4 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ _0776_ _0803_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _0517_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5510_ _2394_ _2389_ _2395_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6490_ mod.des.des_dout\[6\] net4 _3080_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _2268_ _2343_ _2348_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4138__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5335__A1 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5372_ mod.registers.r2\[1\] _2304_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _1203_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout129 net132 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3649__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4310__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ mod.registers.r12\[10\] _1110_ _1106_ mod.registers.r10\[10\] _1155_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__A3 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__B1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3821__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3821__B2 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6698__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _0330_ net46 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4377__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ _0261_ net71 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3969_ _3233_ _0926_ _3249_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5708_ _2528_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _0192_ net57 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5639_ _2472_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3888__B2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A2 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4065__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__B2 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A1 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3812__B2 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4907__A4 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3576__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5317__A1 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3879__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout196_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6045__A2 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4056__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _1909_ _1578_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4851__I0 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6272__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4872_ _1824_ _1836_ _0616_ _0951_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6611_ _0115_ net146 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6990__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ mod.registers.r6\[15\] _0733_ _0766_ mod.registers.r12\[15\] _0793_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3406__I1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3567__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ mod.registers.r15\[13\] _3113_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3754_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5308__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6473_ _2966_ _3044_ _3066_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3685_ mod.registers.r4\[3\] _0508_ _0421_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5859__A2 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ mod.registers.r3\[4\] _2338_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5355_ _2270_ _2290_ _2291_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _1259_ _1271_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5286_ _2201_ _2229_ _2230_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6284__A2 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4237_ _0956_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ mod.registers.r15\[8\] _0963_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4047__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4099_ _1067_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5244__B1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3739__C _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _0313_ net49 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4430__I _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6713__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6863__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__B2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3549__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4340__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3470_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout209_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3316__A3 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5140_ _2094_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6267__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5069__A3 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _2033_ _1963_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4022_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A1 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__B2 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5973_ mod.registers.r14\[13\] _2701_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4924_ _1388_ _1787_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4855_ mod.ldr_hzd\[4\] _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3806_ _0756_ _0775_ _0496_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _1749_ _1753_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6736__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _2410_ _3100_ _3104_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3737_ mod.registers.r11\[3\] _0705_ _0706_ mod.registers.r8\[3\] _0707_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5346__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _2992_ _3061_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3668_ _0637_ _0633_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5407_ _2296_ _2321_ _2326_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4504__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _0862_ _3009_ _3014_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6886__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3599_ mod.registers.r4\[4\] _0420_ _0449_ mod.registers.r1\[4\] _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5338_ _2178_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5269_ _1078_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ _0106_ net205 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4853__C _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3779__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__I0 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6193__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4259__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3482__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4335__I _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout159_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4640_ _0809_ _0842_ _0876_ _0725_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _1241_ _1338_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5931__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5166__I _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6310_ _2961_ _2964_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3522_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ mod.des.des_dout\[7\] _2909_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3453_ _3280_ _3288_ _0414_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6172_ _2753_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3384_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _2056_ _2074_ _2080_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3414__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5054_ _2017_ _1963_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _3178_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3473__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6411__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2410_ _2688_ _2692_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4907_ _1802_ _1810_ _1804_ _1807_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5887_ mod.registers.r12\[13\] _2647_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4973__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4838_ _0637_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4725__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _1280_ _1652_ _1651_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6508_ _3091_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _3048_ _3049_ _3046_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4489__B2 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5150__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4110__B1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__C2 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3464__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6901__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3994__I _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5913__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__B1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__C2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4774__B _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _0294_ net95 mod.registers.r12\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4404__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__B2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ mod.registers.r9\[9\] _2552_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ mod.registers.r8\[3\] _2504_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6213__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4623_ _1409_ _1592_ _1344_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4707__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5904__A1 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3409__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3915__B1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4554_ _1344_ _1356_ _1364_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3915__C2 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3505_ mod.registers.r11\[1\] _3202_ _3195_ mod.registers.r10\[1\] _0475_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4485_ _1097_ _1049_ _1249_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_104_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6224_ _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout91_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5132__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3436_ mod.instr_2\[11\] _3276_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _2833_ _2838_ _2841_ _2847_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ _3212_ _3213_ _3214_ _3218_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5106_ mod.pc0\[9\] _1891_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4684__B _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1943_ _2784_ _1959_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_58_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3298_ mod.des.des_counter\[0\] _3150_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _1998_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6396__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__A2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _0086_ net210 mod.des.des_dout\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3749__A3 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _2679_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6190__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4159__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4174__A3 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3382__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5534__I _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3685__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_225 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3989__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_236 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_247 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_258 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_269 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4398__B1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__B1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4270_ _1004_ _1238_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6947__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__B2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _0009_ net142 mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _0343_ net155 mod.pc0\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3848__B _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ _0277_ net72 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3985_ mod.funct7\[2\] _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5050__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5724_ mod.registers.r9\[4\] _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3600__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5655_ mod.registers.r7\[14\] _2493_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _1366_ _1573_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ _2445_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4537_ _1506_ _1349_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4398__C _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _1253_ _1099_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__B2 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6207_ mod.instr\[0\] _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3419_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4399_ _0934_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6138_ _1913_ _2083_ _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6069_ _1926_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4616__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5529__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6541__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A3 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4589__B _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5264__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3940__C _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3830__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout141_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _0731_ _0734_ _0737_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_20_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5440_ mod.registers.r3\[11\] _2344_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6532__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5335__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5371_ _2177_ _2302_ _2305_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4322_ _1291_ _1220_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5099__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout108 net119 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4253_ _1221_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout119 net128 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3649__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4310__A3 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4184_ mod.registers.r5\[10\] _0882_ _0696_ mod.registers.r4\[10\] _0706_ mod.registers.r8\[10\]
+ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_79_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__B2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3821__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _0329_ net46 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5023__A1 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6756_ _0260_ net140 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3968_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3585__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5707_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6687_ _0191_ net99 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3899_ mod.registers.r13\[9\] _0541_ _0542_ mod.registers.r1\[9\] _0869_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5638_ _2414_ _2480_ _2485_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6523__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5569_ _2295_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3576__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3576__B2 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3879__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4828__A1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout189_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _3243_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3398__B mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__I1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4871_ _1839_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _0114_ net139 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3822_ mod.registers.r5\[15\] _0440_ _0442_ mod.registers.r7\[15\] _0792_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3567__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _2430_ _3112_ _3114_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3753_ _0719_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3567__B2 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _1820_ _3064_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5308__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3684_ mod.registers.r11\[3\] _0505_ _0506_ mod.registers.r2\[3\] _0654_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _2331_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5354_ mod.registers.r1\[14\] _2277_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _1127_ _1150_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ mod.registers.r1\[6\] _2206_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4819__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4236_ _1044_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6665__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4167_ _1135_ _1136_ mod.registers.r1\[8\] _1015_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ _0759_ _0494_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_82_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5244__A1 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5795__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6808_ _0312_ net64 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6739_ _0243_ net125 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__C _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6574__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3997__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5235__A1 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__B2 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3549__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3549__B2 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4210__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout104_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__I _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ mod.pc\[7\] _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__A1 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ _0988_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5972_ _2430_ _2700_ _2702_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6216__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ mod.pc\[0\] _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4017__B _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ mod.ldr_hzd\[5\] _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ _0757_ _0773_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4785_ _1167_ _1669_ _1754_ _1659_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3736_ _3204_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6524_ mod.registers.r15\[6\] _3101_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3667_ _0425_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6455_ _1804_ _3058_ _3059_ _3036_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ mod.registers.r2\[15\] _2322_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6386_ mod.pc_1\[9\] _3010_ _3012_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4687__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3598_ mod.registers.r10\[4\] _3279_ _0413_ mod.registers.r2\[4\] _0568_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3712__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5337_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5268_ _2172_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6501__I1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ _1185_ _1188_ _1181_ _1165_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ _0105_ net204 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _2146_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6407__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3610__I mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4440__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6568__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__I _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6142__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6830__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4597__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3703__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4900__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__I _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5208__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3520__I mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4195__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _0989_ _1538_ _1422_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _0490_ _0482_ _3258_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6479__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _2718_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ mod.registers.r4\[0\] _0420_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6171_ _2781_ _2859_ _2863_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3383_ _3234_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5122_ _2005_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ mod.pc\[6\] _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5998__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4004_ _0605_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3430__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5955_ mod.registers.r14\[6\] _2689_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _1831_ _1847_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5886_ _2560_ _2646_ _2648_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4837_ mod.ldr_hzd\[8\] _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4261__I _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6853__CLK net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _1281_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5922__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6507_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3719_ _0470_ _0488_ _0560_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4699_ _0945_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _2967_ _1862_ _3038_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4489__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__A1 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6369_ _0651_ _3000_ _3002_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__A1 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__B2 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6137__B mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4661__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3340__I mod.instr_2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3621__B1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5267__I _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__A1 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3924__B2 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5677__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5429__A1 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4101__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout171_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3860__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4404__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6876__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ _2253_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__B1 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6157__A2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _2397_ _2502_ _2507_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4168__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4622_ _0529_ _0773_ _0681_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3915__A1 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4553_ _1383_ _1513_ _1516_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3915__B2 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3504_ mod.registers.r8\[1\] _0473_ _3199_ mod.registers.r9\[1\] _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4484_ _1269_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5668__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _2717_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3435_ mod.registers.r14\[0\] _3283_ _3287_ mod.registers.r6\[0\] _3288_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _2774_ _2848_ _2849_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout84_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3366_ mod.registers.r15\[0\] _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ mod.pc\[9\] _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6085_ _2768_ _2769_ mod.pc\[3\] _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5640__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3297_ _3152_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ mod.pc0\[5\] _1960_ _1961_ _2000_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4643__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3851__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _0085_ net210 mod.des.des_dout\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6396__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6404__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ mod.registers.r12\[6\] _2635_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4159__B2 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3906__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3382__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 net23 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_226 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6084__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_237 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_248 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_259 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5831__A1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6899__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6387__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__B2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5898__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5822__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _0008_ net169 mod.instr_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6841_ _0342_ net156 mod.pc0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4389__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6772_ _0276_ net135 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5050__A2 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5723_ _2531_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5654_ _2436_ _2492_ _2495_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5889__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _1555_ _1349_ _1371_ _1450_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5585_ _2400_ _2446_ _2452_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4561__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4536_ _1148_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _1097_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6302__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _2131_ _2883_ _2886_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3418_ _3267_ _3269_ _3270_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4398_ _1362_ _1363_ _1365_ _0627_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _2802_ _1885_ mod.pc\[10\] _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3349_ _3201_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _1911_ _2004_ _1920_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_58_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4077__B1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ _3153_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A3 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6376__I _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__B1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A1 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3815__B1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3949__B _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5032__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4240__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout134_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5370_ mod.registers.r2\[0\] _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4321_ mod.pc_2\[12\] _1205_ _1289_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_126_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5099__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__A1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _0755_ _1220_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ mod.registers.r15\[10\] _0884_ _0879_ mod.registers.r7\[10\] mod.registers.r3\[10\]
+ _0694_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_80_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5190__I _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4059__B1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__C _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5271__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout47_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _0328_ net54 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _0259_ net138 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3967_ _0931_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5706_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6686_ _0190_ net102 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ mod.registers.r15\[9\] _0435_ _0437_ mod.registers.r12\[9\] _0868_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5637_ mod.registers.r7\[7\] _2481_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4534__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3337__A2 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _2439_ _2432_ _2440_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4519_ _1462_ _1465_ _1466_ _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_104_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5499_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6287__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3648__I0 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__C _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3769__B _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__B1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3576__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5275__I _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__B _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4828__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A2 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__I2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4870_ _1815_ _1834_ _1836_ _1813_ _1812_ _1832_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_32_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3821_ mod.registers.r13\[15\] _0745_ _0732_ mod.registers.r14\[15\] _0791_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6540_ mod.registers.r15\[12\] _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4764__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3567__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3752_ _3239_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _3070_ _3071_ _3057_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3683_ mod.registers.r14\[3\] _0534_ _0535_ mod.registers.r6\[3\] _0653_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6505__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3319__A2 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _2329_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4304_ _1272_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5284_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4235_ _0778_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5492__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _0483_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4097_ mod.pc_2\[1\] _0777_ _1065_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6441__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5244__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__A3 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6807_ _0311_ net64 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4055__I0 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1959_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4755__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _0242_ net126 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _0173_ net98 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3608__I _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4507__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5235__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6590__S _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3549__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net82 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net94 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ _0989_ _0986_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4793__B _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ mod.registers.r14\[12\] _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4985__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4853_ _1822_ _1809_ _0636_ _0424_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3804_ _0552_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4784_ _1400_ _1595_ _1481_ _1317_ _1660_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _2407_ _3100_ _3103_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3735_ _3202_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4033__B _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6454_ _2992_ _3060_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3666_ _0562_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _2290_ _2321_ _2325_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _0843_ _3009_ _3013_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6632__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3597_ _0558_ _0559_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3712__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5336_ mod.des.des_dout\[33\] _2248_ _2272_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _2165_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7006_ _0104_ net204 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4218_ _1186_ _1187_ _1126_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5198_ _2147_ _2143_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ mod.registers.r15\[9\] _0884_ _0600_ mod.registers.r6\[9\] _0473_ mod.registers.r8\[9\]
+ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_56_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3779__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__C1 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3338__I _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3703__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6585__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6405__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__B _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3957__B _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4195__A2 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3520_ mod.instr_2\[4\] _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5144__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3451_ _3236_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6170_ mod.pc_1\[1\] _2861_ _2822_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3382_ _3230_ _3231_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4079__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5121_ _2060_ _2078_ _2076_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6495__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5447__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ _1911_ _2004_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A3 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4003_ mod.registers.r4\[15\] _0971_ _0972_ mod.registers.r10\[15\] _0973_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3711__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__B2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _2407_ _2688_ _2691_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__C _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4905_ _1831_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5885_ mod.registers.r12\[12\] _2647_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4836_ _3275_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5383__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _1728_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6506_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3718_ _0687_ _0492_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _1665_ _1666_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6437_ _1825_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3649_ _0615_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6368_ mod.pc_1\[3\] _3001_ _2996_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3697__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4894__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ mod.des.des_dout\[31\] _2248_ _2257_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _0905_ _2956_ _2951_ mod.instr\[0\] _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6486__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3621__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3621__B2 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4177__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5126__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3688__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4885__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3860__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3860__B2 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__B2 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4362__I _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ mod.registers.r8\[2\] _2504_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4621_ _0827_ _0841_ _0802_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4168__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4552_ _1520_ _1521_ _1432_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3915__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _3203_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4483_ _1449_ _1451_ _1452_ _1445_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5193__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ mod.instr\[3\] _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3434_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ mod.pc\[12\] _2774_ _2822_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3365_ _3215_ _3216_ _3209_ _3217_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _2056_ _2055_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout77_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _1944_ _2780_ _2787_ _2789_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3296_ net165 _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _1999_ _1963_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4643__A3 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__A1 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3851__B2 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _0084_ net212 mod.des.des_dout\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3603__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4272__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ _2544_ _2634_ _2637_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5356__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4159__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _0902_ _1785_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6970__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5799_ _2560_ _2591_ _2593_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3367__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3906__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput24 net24 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4867__B1 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4867__C2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_227 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_238 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_249 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3351__I _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5831__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4182__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3526__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4357__I _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6843__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3833__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6840_ _0341_ net156 mod.pc0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6993__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6771_ _0275_ net135 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3983_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5188__I _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ _2529_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ mod.registers.r7\[13\] _2493_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5916__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _1068_ _0933_ _0939_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5584_ mod.registers.r6\[3\] _2448_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4535_ _1327_ _0810_ _0877_ _1339_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4466_ _1242_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6205_ mod.pc_1\[13\] _2884_ _2880_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4313__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5510__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3417_ mod.instr_2\[11\] mod.instr_2\[10\] _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4397_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _2833_ _2829_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3348_ _3196_ _3197_ _3160_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4077__B2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5018_ _1969_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _0067_ net214 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3588__B1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5329__A1 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6716__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3346__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5561__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4068__B2 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3815__A1 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3815__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4083__A4 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4240__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4240__B2 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4791__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5736__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout127_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _0742_ _0744_ _0750_ _0753_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__3897__A4 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__B _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6567__I _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4251_ _0755_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4182_ _0489_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6048__A2 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4059__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4059__B2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3806__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6823_ _0327_ net53 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6754_ _0258_ net138 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3966_ _3226_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4231__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4231__B2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6739__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5705_ _2161_ _2499_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4782__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6685_ _0189_ net98 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3897_ _0863_ _0864_ _0865_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5636_ _2411_ _2480_ _2484_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5731__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ mod.registers.r5\[14\] _2433_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3337__A3 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6889__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ _1224_ _1397_ _1479_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _2176_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__A2 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _0715_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6119_ _2033_ _2780_ _2819_ _2789_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5798__A1 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3648__I1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4470__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6598__I0 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4222__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__B2 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__I _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A2 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4851__I3 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3820_ _0779_ _0789_ _0556_ _0557_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3751_ _0720_ _0712_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4764__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5961__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4370__I _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _3055_ _3041_ _3066_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3682_ mod.registers.r8\[3\] _0531_ _0532_ mod.registers.r10\[3\] _0652_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5421_ _2199_ _2330_ _2336_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4516__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ mod.des.des_dout\[35\] _2220_ _2286_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_114_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4303_ _1180_ _1181_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6297__I _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5283_ mod.des.des_dout\[27\] _2220_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3714__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4234_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4165_ _3183_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _0675_ _0676_ _0677_ _0678_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4452__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6806_ _0310_ net69 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4204__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ mod.pc0\[3\] _1960_ _1961_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4055__I1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6737_ _0241_ net126 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3949_ _0718_ _0913_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5952__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6668_ _0172_ net85 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ _2471_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6599_ _3147_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__I _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6904__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout70 net73 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout81 net83 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3706__B1 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5235__B _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout194_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3485__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _2682_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4985__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6580__I _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ mod.ldr_hzd\[6\] _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6187__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3803_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4198__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__C2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5934__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _1750_ _1751_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6522_ mod.registers.r15\[5\] _3101_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ mod.registers.r10\[3\] _0602_ _0703_ mod.registers.r9\[3\] _0704_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _1807_ _3058_ _3059_ _1862_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3665_ _0631_ _0632_ mod.registers.r11\[2\] _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5404_ mod.registers.r2\[14\] _2322_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6384_ mod.pc_1\[8\] _3010_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3596_ mod.registers.r13\[4\] _0447_ _0431_ mod.registers.r3\[4\] _0565_ _0566_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5335_ _2025_ _2273_ _2166_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3712__A3 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6111__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _0580_ _2189_ _2209_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6927__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7005_ _0103_ net219 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4217_ _0859_ _1147_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5197_ mod.rd_3\[3\] _2144_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3476__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _1114_ _1115_ _1116_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_83_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6414__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3779__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4728__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__C2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4113__B1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4195__A3 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout207_I net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3381_ mod.instr_2\[1\] _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5120_ _2077_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ _2005_ _2007_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4002_ _0602_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ mod.registers.r14\[5\] _2689_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5080__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1866_ _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5884_ _2628_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4835_ _0633_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3439__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _1332_ _1731_ _1732_ _1735_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3717_ _0615_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6505_ _2327_ _2624_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4697_ _1307_ _1544_ _0922_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ _3032_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3648_ mod.instr_2\[5\] _0616_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6367_ _2952_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3579_ mod.registers.r5\[7\] _0547_ _0548_ mod.registers.r7\[7\] _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3697__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__B2 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ _2174_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6298_ _2955_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _0651_ _2168_ _2173_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4646__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4219__B _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5829__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3621__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3349__I _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3793__B _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6596__S _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3688__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4885__B2 mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4637__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3860__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout157_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6622__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3612__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _1267_ _1349_ _0921_ _1587_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5365__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1438_ _1519_ _1495_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3502_ mod.registers.r3\[1\] _0471_ _3186_ mod.registers.r6\[1\] mod.registers.r7\[1\]
+ _3170_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_4482_ _1056_ _1061_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6221_ _2895_ _2719_ _2897_ _2892_ _2898_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3433_ _3284_ _3285_ _3274_ _3276_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _2845_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _3159_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _2059_ _2062_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6083_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3295_ _0000_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ mod.pc\[5\] _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3300__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4643__A4 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3851__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _0083_ net48 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5649__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _2299_ _2624_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4800__A1 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3603__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ mod.registers.r12\[5\] _2635_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5356__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5798_ mod.registers.r10\[12\] _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4749_ _1713_ _1714_ _1715_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_31_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5108__A2 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput25 net25 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _1812_ _0003_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_89_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput36 net36 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4867__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4867__B2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3632__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6148__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_228 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_239 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3827__C1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4634__A4 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6645__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4463__I _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6795__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6544__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3542__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__S _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3833__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4373__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3982_ _3232_ _3252_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6770_ _0274_ net134 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ _2204_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _2431_ _2492_ _2494_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4603_ _1309_ _1333_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5583_ _2397_ _2446_ _2451_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3717__I _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4534_ _1420_ _1502_ _1503_ _0920_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6299__B1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4465_ _1398_ _1428_ _1431_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_3416_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6204_ _2115_ _2883_ _2885_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4396_ _0725_ _0920_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4548__I _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6135_ _2816_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3347_ mod.registers.r10\[0\] _3195_ _3199_ mod.registers.r9\[0\] _3200_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6668__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _2726_ _1900_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5017_ _1979_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5379__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4283__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6968_ _0066_ net211 mod.des.des_dout\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3588__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3588__B2 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__B1 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5919_ _2416_ _2667_ _2669_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6899_ _0400_ net165 mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__I _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__I1 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6159__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3815__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3579__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3579__B2 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4240__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _1205_ _1208_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4059__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6453__B1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6822_ _0326_ net60 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _0257_ net138 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5927__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3965_ mod.funct3\[0\] _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4231__A2 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5704_ _2176_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6684_ _0188_ net41 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3896_ mod.registers.r4\[9\] _0508_ _0421_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ mod.registers.r7\[6\] _2481_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5566_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4517_ _1332_ _1483_ _1486_ _1222_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5497_ _2296_ _2379_ _2384_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5662__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4448_ _1400_ _1408_ _1417_ _1329_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5495__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4379_ _3229_ _3244_ _3247_ _0936_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _2814_ _2817_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ _2741_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6598__I1 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6442__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4222__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6161__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6833__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6983__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5486__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3497__B1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3976__B _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3750_ _0560_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5961__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3681_ mod.pc_2\[3\] _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5420_ mod.registers.r3\[3\] _2332_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _2220_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4302_ _1165_ _1166_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5282_ _2222_ _2223_ _2225_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4233_ _0772_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _0711_ _1113_ mod.registers.r8\[8\] _1010_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5229__A1 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3730__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _0670_ _0671_ _0672_ _0673_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout52_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6805_ _0309_ net69 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5401__A1 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4997_ _1962_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4204__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6856__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _0240_ net70 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3948_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__A3 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6667_ _0171_ net84 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3879_ mod.registers.r12\[8\] _0848_ _0638_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5618_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6598_ net6 mod.des.des_dout\[34\] _3136_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5549_ mod.registers.r5\[10\] _2419_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout60 net61 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout71 net73 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A1 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3706__B2 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4131__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3485__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout187_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3550__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6879__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4920_ _1884_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3642__B1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _1817_ _1818_ _1819_ _1820_ _1805_ _1808_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6187__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3802_ _0758_ _0759_ _0764_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4198__B2 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5934__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4782_ _1467_ _1587_ _1329_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6521_ _2402_ _3100_ _3102_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3733_ _3198_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _2147_ _2966_ _3025_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3664_ _0444_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5698__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2284_ _2321_ _2324_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3595_ _0560_ _0561_ _0563_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6383_ _2752_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5334_ _2224_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _2210_ _1988_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5940__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4122__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7004_ _0102_ net204 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4216_ _0874_ _1124_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5196_ _1848_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5870__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4673__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3476__A3 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4147_ _0951_ _0616_ mod.registers.r4\[9\] _1010_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ _0524_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4505__B _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4189__B2 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _0223_ net100 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5689__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__I _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4113__B2 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3370__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5613__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3545__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout102_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5760__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1790_ _2013_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ _3174_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5604__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _2402_ _2688_ _2690_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ mod.instr_2\[6\] _1869_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _2626_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4834_ mod.ldr_hzd\[9\] _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _1204_ _1397_ _1546_ _1330_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _3090_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3716_ _0682_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _1322_ _1355_ _0497_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _3043_ _3045_ _3046_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4060__B _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3647_ _3258_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6366_ _2713_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3578_ _0441_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4894__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1991_ _2226_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _2856_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6096__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _2169_ _1950_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5843__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5179_ _2072_ _2120_ _2134_ _3156_ _2135_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4219__C _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6020__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4582__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4885__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A1 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3845__B1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6917__CLK net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4550_ _1438_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3501_ _3164_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _1068_ _1450_ _0454_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6220_ _2788_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3432_ mod.instr_2\[12\] _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _2114_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3363_ _3162_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _2059_ _2062_ _1790_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _2706_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3294_ mod.des.des_counter\[1\] _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _1934_ _1912_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_38_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3300__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _0082_ net47 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6254__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ _2441_ _2673_ _2678_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5866_ _2540_ _2634_ _2636_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6002__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0908_ _1784_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_21_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ _2573_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5356__A3 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5665__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4564__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3367__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _1716_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _1259_ _1271_ _1492_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6418_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput26 net26 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput37 net37 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6349_ _0711_ _2989_ _2986_ mod.instr\[17\] _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5816__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_229 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3827__B1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3827__C2 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4095__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5575__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5283__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _3196_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5720_ _2538_ _2530_ _2539_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ mod.registers.r7\[12\] _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6090__B _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6535__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ _1382_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5582_ mod.registers.r6\[2\] _2448_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _0924_ _0927_ _0717_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6299__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6299__B2 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _1302_ _1296_ _1399_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_89_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6203_ mod.pc_1\[12\] _2884_ _2880_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3415_ mod.instr_2\[12\] _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4395_ _1226_ _1357_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3733__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout82_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6134_ mod.pc\[10\] _2824_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _1893_ _2766_ _2772_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5274__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ mod.pc0\[4\] _1922_ _1923_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _0065_ net211 mod.des.des_dout\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4785__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ mod.registers.r13\[8\] _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3588__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4785__B2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6898_ _0399_ net165 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ _2355_ _2498_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3908__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4513__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6762__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3579__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4423__B _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3751__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _1148_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6453__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__B2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5008__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6821_ _0325_ net61 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _0256_ net71 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3964_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ _2442_ _2521_ _2526_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4231__A3 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6683_ _0187_ net41 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3895_ mod.registers.r11\[9\] _3292_ _0506_ mod.registers.r2\[9\] _0865_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5148__C _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _2408_ _2480_ _2483_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5565_ _2289_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ _1228_ _1369_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ mod.registers.r4\[15\] _2380_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4447_ _1400_ _1412_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3463__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4378_ _1332_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _2764_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ mod.instr_2\[15\] _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6444__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _2730_ _2105_ _2758_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3373__I mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3497__A1 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5238__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__A3 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3548__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3680_ _0628_ _0577_ _0643_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _1233_ _2273_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _1263_ _1268_ _1269_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_5_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _2171_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4232_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ mod.registers.r6\[8\] _0700_ _0696_ mod.registers.r4\[8\] _0603_ mod.registers.r9\[8\]
+ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4328__B _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4094_ _1055_ _1061_ _1062_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_55_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4988__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5003__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout45_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5938__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3660__B2 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6804_ _0308_ net116 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6262__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4996_ _1924_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5401__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _0239_ net109 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3947_ _3227_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3458__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _0170_ net85 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3878_ _0631_ _0562_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5165__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6597_ _3146_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4912__A1 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4912__B2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6114__B1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5479_ _2361_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3921__I _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6417__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4691__A3 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6800__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout72 net73 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout83 net86 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3954__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3706__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__B1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3831__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5631__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6363__B _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3642__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3642__B2 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ mod.ldr_hzd\[15\] _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3801_ _0767_ _0768_ _0769_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4198__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5395__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _1352_ _1404_ _1473_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ mod.registers.r15\[4\] _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3732_ mod.registers.r6\[3\] _0700_ _0468_ mod.registers.r5\[3\] mod.registers.r2\[3\]
+ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5147__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _3032_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _3276_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ mod.registers.r2\[13\] _2322_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6382_ _0530_ _3009_ _3011_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3594_ mod.registers.r15\[4\] _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _2123_ _2189_ _2214_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5264_ _1793_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _0101_ net208 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4215_ _1166_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4837__I mod.ldr_hzd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3741__I _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _2141_ _2143_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4146_ _0482_ _0483_ mod.registers.r13\[9\] _0478_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3881__A1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6823__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4077_ _1021_ _1043_ _1046_ _0458_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_71_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4505__C _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A1 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4979_ _1943_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6718_ _0222_ net100 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _0153_ net80 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__B1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__A2 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5613__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4352__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4104__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5301__A1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3561__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6846__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ _0961_ _0965_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5951_ mod.registers.r14\[4\] _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6093__B mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6996__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _1870_ _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5882_ _2558_ _2640_ _2645_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _1802_ _0429_ _0632_ _0846_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _0922_ _1733_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6503_ mod.des.des_dout\[12\] net10 _3074_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3715_ _0683_ _0684_ _0453_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4695_ _1315_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3736__I _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6434_ _2715_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5156__C _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3646_ _3216_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _0628_ _2714_ _2999_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3577_ _0439_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _2075_ _2189_ _2209_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2951_ _2954_ _2831_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5247_ _2164_ _2194_ _2195_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _3154_ _2122_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _1093_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4516__B _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5398__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5359__A1 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4031__A1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4582__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6869__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3381__I mod.instr_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3845__A1 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3845__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5598__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5257__B _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3556__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout212_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3500_ _0467_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4480_ _0688_ _0689_ _1069_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3431_ mod.instr_2\[13\] _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6570__I0 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3679__A4 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ mod.pc\[12\] _1914_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _3181_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _2060_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4387__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _2765_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3293_ mod.des.des_counter\[0\] _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__B2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _1915_ _1988_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5038__B1 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5589__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6983_ _0081_ net46 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ mod.registers.r13\[15\] _2674_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ mod.registers.r12\[4\] _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6002__A2 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4816_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ _2571_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5356__A4 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _1030_ _1669_ _1485_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4564__A2 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4678_ _1280_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6417_ _2728_ _1801_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3629_ _0597_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5513__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput27 net27 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput38 net38 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6348_ _2860_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ mod.instr\[17\] _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3827__B2 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6017__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5752__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6691__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout162_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3980_ _0779_ _0878_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5650_ _2474_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4601_ _1563_ _1567_ _1570_ _0918_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5581_ _2394_ _2446_ _2450_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4532_ _1500_ _1470_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4463_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6202_ _2857_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3414_ mod.instr_2\[13\] _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4394_ _0529_ _1291_ _0553_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_112_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _2825_ _2830_ _2831_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3345_ _3196_ _3197_ _3175_ _3187_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _2767_ _2771_ _2754_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout75_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _1980_ _1897_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6265__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6966_ _0064_ net214 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _2655_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6897_ _0398_ net184 mod.valid2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _2568_ _2618_ _2623_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5734__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _2540_ _2579_ _2581_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4473__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__A1 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5725__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6150__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _0324_ net123 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4216__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4767__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3963_ _0930_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6751_ _0255_ net111 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ mod.registers.r8\[15\] _2522_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6682_ _0186_ net41 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3894_ mod.registers.r14\[9\] _0534_ _0535_ mod.registers.r6\[9\] _0864_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5716__A1 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ mod.registers.r7\[5\] _2481_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5564_ _2436_ _2432_ _2437_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4515_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _2290_ _2379_ _2383_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _1351_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _1328_ _1335_ _1340_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3328_ _3161_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6047_ _2729_ mod.pc0\[11\] _2754_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4455__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__A2 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _0047_ net174 mod.ldr_hzd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4524__B _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3919__I _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__I _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3497__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout125_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3564__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4300_ _1033_ _1048_ _1094_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5280_ _1046_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4231_ _1135_ _1191_ _0561_ _0985_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ mod.registers.r10\[8\] _1106_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ _0719_ _0722_ _0666_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4988__A2 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3660__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6803_ _0307_ net122 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ mod.pc\[3\] _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6734_ _0238_ net110 mod.registers.r9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3946_ _0914_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6665_ _0169_ net85 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3877_ _0846_ _0632_ mod.registers.r11\[8\] _0634_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5616_ _2327_ _2356_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5165__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ net5 mod.des.des_dout\[33\] _3142_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6752__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _2260_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6114__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _2359_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4429_ _1237_ _1287_ _1295_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_78_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4676__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5928__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6025__I _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout40 net42 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout51 net52 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4600__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout62 net63 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout73 net74 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout84 net86 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5864__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3384__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6105__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4116__B1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4667__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6408__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4943__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6625__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3642__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3559__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ mod.registers.r5\[13\] _0741_ _0743_ mod.registers.r7\[13\] _0770_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4780_ _1665_ _1415_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3731_ _3190_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3945__A3 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6450_ _3054_ _3056_ _3057_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6344__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3662_ _0416_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6344__B2 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5401_ _2276_ _2321_ _2323_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6381_ mod.pc_1\[7\] _3010_ _3004_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3593_ _0415_ _0562_ _0444_ _3277_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_127_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5332_ _2210_ _2108_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4214_ _1102_ _1105_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7002_ _0100_ net205 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5194_ mod.rd_3\[2\] _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4145_ _0480_ _3256_ mod.registers.r14\[9\] _0478_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5014__I mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _1044_ _0491_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ mod.pc0\[2\] _1922_ _1923_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3397__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6717_ _0221_ net109 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3929_ _0759_ _0896_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5684__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _0152_ net87 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6335__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6335__B2 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3932__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__B2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6648__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3872__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4121__I0 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3624__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4821__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6798__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3388__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5129__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout192_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _2682_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4812__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3615__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ mod.ldr_hzd\[8\] _1856_ _1858_ mod.ldr_hzd\[10\] mod.instr_2\[5\] _1871_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ mod.registers.r12\[11\] _2641_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4832_ mod.ldr_hzd\[11\] _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3379__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4763_ _1333_ _1365_ _0627_ _1359_ _1666_ _1343_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _3089_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3714_ _0557_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4694_ _1659_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _3029_ _3044_ _3038_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3645_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6364_ mod.pc_1\[2\] _2995_ _2996_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3576_ mod.registers.r9\[7\] _0544_ _0545_ mod.registers.r3\[7\] _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5315_ _2210_ _2074_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6295_ _1886_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5246_ mod.registers.r1\[2\] _2179_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ _2130_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _1076_ _1093_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5056__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4059_ mod.pc_2\[7\] _0499_ _1027_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5359__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4031__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__A1 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3790__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A1 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout205_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6369__B _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6570__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3361_ _3206_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3572__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ mod.pc_2\[9\] _1233_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _2783_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6963__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _1916_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5038__A1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5499__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _0080_ net47 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5589__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _2438_ _2673_ _2677_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4797__B1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _2628_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _0904_ _0905_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3747__I _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ _2558_ _2585_ _2590_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4746_ _1031_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5761__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3772__A1 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _1511_ _1554_ _1579_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ _2147_ _2956_ _3031_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3628_ mod.registers.r4\[2\] _3174_ _3178_ mod.registers.r1\[2\] _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6561__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput28 net28 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6347_ _2985_ _2988_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3559_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6278_ _2939_ _2937_ _2940_ _2941_ _2935_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5277__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ mod.registers.r1\[0\] _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3827__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5201__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5752__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__A3 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6552__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6986__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3392__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__C1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__B1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout155_I net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _0726_ _1568_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4546__A3 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ mod.registers.r6\[1\] _2448_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _1305_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4462_ _3250_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ _2867_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3413_ _3265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4393_ _0925_ _1334_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _2707_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3344_ mod.instr_2\[16\] _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _1797_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ mod.pc\[4\] _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout68_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5022__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _0063_ net214 mod.des.des_dout\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5431__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5916_ _2653_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _0397_ net170 mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5847_ mod.registers.r11\[15\] _2619_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3477__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5778_ mod.registers.r10\[4\] _2580_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3745__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _1429_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4170__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5670__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4225__A2 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4704__C _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4011__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5110__B1 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5661__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__B _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5777__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4216__A2 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _0254_ net111 mod.registers.r10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3962_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5701_ _2439_ _2521_ _2525_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6681_ _0185_ net41 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3893_ mod.registers.r8\[9\] _3273_ _0532_ mod.registers.r10\[9\] _0863_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6602__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5632_ _2403_ _2480_ _2482_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5563_ mod.registers.r5\[13\] _2433_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6401__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4514_ _0937_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5494_ mod.registers.r4\[14\] _2380_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4445_ _1413_ _1414_ _1313_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _1343_ _1345_ _1336_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _2782_ _2791_ _2807_ _2815_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3327_ _3171_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2743_ _2757_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6681__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A1 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _0046_ net177 mod.ldr_hzd\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3966__A1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _0380_ net176 mod.instr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3935__I _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__A3 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5891__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4446__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__A1 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3957__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ _1152_ _1196_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4685__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4161_ _1129_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3893__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _3245_ _0714_ _1059_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_370 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _0306_ net124 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4994_ _1899_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6733_ _0237_ net109 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3945_ _3228_ _3233_ _0728_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4070__B1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6664_ _0168_ net88 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3876_ _0631_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _2442_ _2465_ _2470_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3755__I _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6362__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _3145_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5546_ _2422_ _2418_ _2423_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5477_ _2236_ _2367_ _2372_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5970__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4125__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4428_ _1396_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4676__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4359_ _0920_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3884__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__C _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4428__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5625__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _2743_ _2745_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3636__B1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4535__B _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6306__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout41 net43 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4600__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net76 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout63 net75 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout96 net97 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6041__I _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4364__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4116__B2 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3614__B _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3875__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5616__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3627__B1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5092__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3730_ _3185_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3575__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3661_ _0415_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4355__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ mod.registers.r2\[12\] _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6380_ _2952_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3592_ _3268_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _2163_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4107__A1 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _2172_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4658__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7001_ _0099_ net208 mod.des.des_dout\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _1128_ _1151_ _1167_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5193_ _2142_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3866__B1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4144_ _3215_ _1113_ mod.registers.r11\[9\] _1013_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ mod.funct3\[1\] _1024_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3618__B1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout50_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6032__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ _1944_ _1897_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ _0220_ net39 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4594__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3397__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3928_ _0720_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6647_ _0151_ net90 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ mod.registers.r8\[10\] _0729_ _0730_ mod.registers.r10\[10\] _0829_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6335__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ mod.des.des_counter\[2\] _2071_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _2228_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5846__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3872__A3 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5074__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4821__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__A2 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__I _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5837__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__I mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout185_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6262__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6742__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ mod.ldr_hzd\[11\] _1852_ _1854_ mod.ldr_hzd\[9\] _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ _2556_ _2640_ _2644_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ net14 _1798_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4025__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3379__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1227_ _1485_ _1369_ _1229_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4576__B2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ mod.des.des_dout\[11\] net9 _3085_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _0556_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4693_ _1660_ _1661_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4328__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6432_ _1852_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3644_ _0456_ _3235_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _0669_ _2714_ _2998_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3575_ _0430_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5314_ _2238_ _2254_ _2255_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _2952_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5828__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5245_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ mod.pc0\[13\] _1892_ _1901_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__I _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ _1032_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__C _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4058_ _0540_ _0543_ _0546_ _0549_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5695__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4567__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4319__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3790__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6615__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4098__A3 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6765__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6906__D _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6547__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3360_ _3172_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5286__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ mod.pc_2\[5\] _1991_ _1994_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_85_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6385__B _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6981_ _0079_ net65 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4246__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ mod.registers.r13\[14\] _2674_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4797__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _2626_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4633__B _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4549__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _1390_ _1393_ _1777_ _1780_ _1783_ _1391_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5794_ mod.registers.r10\[11\] _2586_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4013__A3 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5210__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _1030_ _1670_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6638__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3772__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4676_ _1604_ _1621_ _1627_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6415_ mod.rd_3\[3\] _2858_ _2140_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3627_ mod.registers.r3\[2\] _3165_ _0596_ mod.registers.r7\[2\] _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3763__I _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput29 net29 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ _0616_ _2982_ _2986_ mod.instr\[16\] _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3524__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3558_ _0464_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ net13 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3489_ _0457_ _3259_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5277__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5159_ mod.pc0\[12\] _1891_ _1900_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4788__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3460__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4712__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__C _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4228__C2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout148_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ _1474_ _1475_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4461_ _1238_ _1429_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3583__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6200_ _2102_ _2876_ _2882_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3412_ _3264_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4392_ _0789_ _0813_ _0814_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _2826_ _2827_ _2829_ _2817_ _2773_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _3193_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2768_ _2769_ mod.pc\[0\] _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _1934_ _1912_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _0062_ net213 mod.des.des_dout\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _2413_ _2661_ _2666_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6895_ _0396_ net170 mod.instr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3758__I _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _2566_ _2618_ _2622_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _2573_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4728_ _1435_ _1489_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_108_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4659_ _1353_ _1525_ _0496_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _1805_ _2975_ _2972_ mod.instr\[10\] _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6803__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__B1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6953__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5661__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3228_ _3240_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3578__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ mod.registers.r8\[14\] _2522_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ _0184_ net55 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3892_ mod.pc_2\[9\] _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5177__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ mod.registers.r7\[4\] _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5562_ _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4924__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4513_ _1473_ _1482_ _1340_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5493_ _2284_ _2379_ _2382_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _1357_ _0840_ _0875_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4375_ _1344_ _0527_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6429__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _2016_ _2809_ _2032_ _2813_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ mod.registers.r4\[0\] _3174_ _3178_ mod.registers.r1\[0\] _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _2746_ mod.pc0\[10\] _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6826__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__C _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A3 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6947_ _0045_ net175 mod.ldr_hzd\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4093__B _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3488__I _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _0379_ net176 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5168__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _2598_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3718__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__I _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5643__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3654__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3957__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__B1 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__B2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6849__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ mod.registers.r14\[8\] _0891_ _0889_ mod.registers.r13\[8\] _1130_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3893__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3893__B2 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _0804_ _0806_ _0650_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_110_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6999__CLK net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_360 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_371 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _0305_ net114 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4993_ _1890_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6732_ _0236_ net39 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3944_ mod.funct3\[0\] _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4070__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4070__B2 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6663_ _0167_ net88 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3875_ mod.registers.r7\[8\] _0442_ _3287_ mod.registers.r6\[8\] _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5614_ mod.registers.r6\[15\] _2466_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ net4 mod.des.des_dout\[32\] _3142_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5545_ mod.registers.r5\[9\] _2419_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ mod.registers.r4\[7\] _2368_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _0945_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4125__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3771__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6287__C _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A3 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__B2 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ mod.instr_2\[16\] _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4289_ _1248_ _1255_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _2734_ mod.pc0\[5\] _2744_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3636__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__B2 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3939__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4061__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout42 net43 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A3 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout53 net56 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__B _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout64 net68 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout75 net76 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout86 net96 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net152 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5313__A1 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4116__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__I mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3875__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3875__B2 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5616__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3627__B2 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3856__I _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout130_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ mod.registers.r14\[2\] _0534_ _0535_ mod.registers.r6\[2\] _0630_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4355__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3591_ _3235_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6671__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _2238_ _2268_ _2269_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3563__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _2201_ _2205_ _2207_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5304__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7000_ _0098_ net208 mod.des.des_dout\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4212_ _1180_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5855__A2 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5192_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3866__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3866__B2 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4143_ _3168_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4074_ _1024_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3618__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3618__B2 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4291__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout43_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4043__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4976_ mod.pc\[2\] _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ _0219_ net43 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4594__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3766__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3397__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5791__A1 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ mod.funct7\[1\] mod.funct7\[0\] _0617_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3858_ _0728_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6646_ _0150_ net87 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6577_ _3134_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3789_ _0458_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5981__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3554__B1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5528_ _2408_ _2404_ _2409_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3715__B _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5459_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_120_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A2 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5782__A1 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5837__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3848__A1 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout178_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ net15 _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4025__A1 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4025__B2 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4761_ _1473_ _1730_ _1340_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4576__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5773__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3586__I _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6500_ _3088_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3712_ _0579_ _0680_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4692_ _1495_ _1338_ _1565_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4328__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3643_ _0601_ _0604_ _0606_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6431_ _1815_ _3033_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6362_ mod.pc_1\[1\] _2995_ _2996_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3574_ _0427_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5313_ mod.registers.r1\[9\] _2246_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6293_ _2712_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5306__I _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5244_ mod.des.des_dout\[23\] _2188_ _2190_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5175_ _2131_ _1925_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _1075_ _1094_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4057_ _0533_ _0536_ _0537_ _0538_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4264__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4880__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4813__C _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _1914_ _1920_ _1927_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _0133_ net92 mod.registers.r2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4120__I mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4255__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4494__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _0078_ net64 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4246__B2 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _2435_ _2673_ _2676_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__A1 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _2538_ _2627_ _2633_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4813_ _1390_ _1776_ _1782_ _0943_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5793_ _2556_ _2585_ _2589_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4744_ _1326_ _1367_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4675_ _1572_ _1623_ _1640_ _1331_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_107_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3626_ _3169_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6414_ _3029_ _2956_ _3030_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6171__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6345_ _2985_ _2987_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3557_ _0460_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3524__A3 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ mod.des.des_dout\[16\] _2933_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _3237_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _2162_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4485__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _2115_ _1925_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4109_ mod.registers.r2\[5\] _3190_ _3169_ mod.registers.r7\[5\] _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _2050_ _1896_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__A1 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6732__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6882__CLK net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4228__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__B2 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5976__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4734__B _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3739__B1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4951__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6240__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _1237_ _1225_ _1230_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__A1 mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3411_ _3236_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4703__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _1352_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5900__A1 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6130_ _2828_ _2827_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3911__B1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3342_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6396__B _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4695__I _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1788_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5012_ _1970_ _1976_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _0061_ net213 mod.des.des_dout\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5967__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6605__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5914_ mod.registers.r13\[7\] _2662_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6894_ _0395_ net145 mod.instr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ mod.registers.r11\[14\] _2619_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ _2571_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6755__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4727_ _1647_ _1674_ _1685_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6144__A1 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _1320_ _1354_ _1406_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3609_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4589_ _1528_ _1529_ _1342_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _2971_ _2976_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4170__A3 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6259_ mod.instr\[12\] _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4458__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4464__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout160_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _3248_ _0914_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4621__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6778__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3891_ _0552_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _2474_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6374__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5561_ _2283_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4924__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3594__I mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4512_ _1307_ _1480_ _1481_ _1337_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6126__A1 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5492_ mod.registers.r4\[13\] _2380_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4137__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _0554_ _0860_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4688__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4374_ _0625_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6113_ _2808_ _2810_ _2032_ _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3325_ _3177_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6429__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _2722_ _2084_ _2087_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout73_I net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _0044_ net178 mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _0378_ net179 mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5984__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _2548_ _2606_ _2611_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5168__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5759_ _2566_ _2561_ _2567_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4679__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5340__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4549__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6920__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__C1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6356__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__B2 mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A2 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__A1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4390__I0 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3893__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _0723_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_350 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_361 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_372 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _0304_ net110 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4992_ _1934_ _1788_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4445__I1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6731_ _0235_ net47 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3943_ _0726_ _0810_ _0877_ _0901_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4070__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6662_ _0166_ net92 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3874_ mod.registers.r4\[8\] _0420_ _0435_ mod.registers.r15\[8\] _0844_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _2439_ _2465_ _2469_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _3144_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5544_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3581__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__B2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5475_ _2229_ _2367_ _2371_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _1237_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5322__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A4 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ _0716_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__I mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3884__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3308_ mod.instr_2\[17\] _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4288_ _1033_ _1256_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6943__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6027_ _2736_ _1998_ _2001_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _0027_ net162 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout43 net52 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout54 net56 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6338__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout65 net68 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6338__B2 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout76 net97 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout87 net95 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6510__A1 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3324__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6329__B2 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5001__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3590_ _3234_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3563__B2 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ mod.registers.r1\[4\] _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _0825_ _1177_ _1179_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5191_ mod.ins_ldr_3 mod.valid_out3 net15 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_96_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3866__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ mod.registers.r2\[9\] _0701_ _3178_ mod.registers.r1\[9\] _0596_ mod.registers.r7\[9\]
+ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073_ _0489_ _1037_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3618__A2 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4291__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _1934_ _1912_ _1942_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6714_ _0218_ net40 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3926_ _3253_ _0886_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4594__A3 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5791__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6645_ _0149_ net88 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3857_ _0813_ _0814_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6576_ mod.des.des_dout\[25\] net10 _3118_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3788_ mod.pc_2\[13\] _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_164_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3554__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__I mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3554__B2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ mod.registers.r5\[5\] _2405_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3782__I _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _2358_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4409_ _0950_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout200 net201 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout211 net212 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5389_ _2303_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5059__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4282__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A2 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3793__A1 mod.registers.r4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4737__B _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5470__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4025__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5222__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4760_ _1665_ _1535_ _1729_ _1422_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3711_ _3261_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4691_ _1420_ _1568_ _1569_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6430_ _3040_ _3042_ _3023_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3642_ mod.registers.r14\[2\] _0607_ _0608_ mod.registers.r13\[2\] _0611_ _0612_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6361_ _3263_ _2714_ _2997_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3573_ mod.registers.r13\[7\] _0541_ _0542_ mod.registers.r1\[7\] _0543_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5312_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6292_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5289__A1 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5243_ _0628_ _2191_ _2174_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ mod.pc\[13\] _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ _0899_ _0574_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6418__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _0458_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4264__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3777__I mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _1921_ _1922_ _1923_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3909_ _3170_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5992__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4889_ mod.ldr_hzd\[0\] _1856_ _1858_ mod.ldr_hzd\[2\] mod.instr_2\[5\] _1859_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6628_ _0132_ net139 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ mod.des.des_dout\[17\] net2 _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6661__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5691__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3371__B _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout190_I net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ mod.registers.r13\[13\] _2674_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5994__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ mod.registers.r12\[3\] _2629_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _1781_ _1394_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5792_ mod.registers.r10\[10\] _2586_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ _1708_ _1711_ _1712_ _1332_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4674_ _1366_ _1641_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3509__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6413_ mod.rd_3\[2\] _2858_ _2140_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3625_ _0489_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6171__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6344_ _0480_ _2982_ _2986_ mod.instr\[15\] _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3556_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6459__B1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6275_ mod.instr\[16\] _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3487_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5226_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__A1 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6684__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ mod.pc\[12\] _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3693__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _1024_ _3259_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ mod.pc\[8\] _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5987__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input16_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4891__I mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ mod.registers.r12\[7\] _0888_ _0608_ mod.registers.r13\[7\] _1009_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4788__A3 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3920__B2 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3739__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__B2 mod.registers.r13\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6153__A2 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3410_ mod.pc_2\[0\] _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__4164__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1355_ _1359_ _0497_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4976__I mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3341_ _3193_ _3162_ _3182_ _3184_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1389_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ _1794_ _1968_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4219__A2 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5416__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _0060_ net213 mod.des.des_dout\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3427__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5967__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3978__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _2410_ _2661_ _2665_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6893_ _0394_ net145 mod.instr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _2564_ _2618_ _2621_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ _2538_ _2572_ _2578_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4726_ _3242_ _1680_ _1691_ _1659_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_108_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _1301_ _1623_ _1626_ _1432_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_107_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4155__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4588_ _1556_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ _1781_ _2975_ _2972_ mod.instr\[9\] _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3539_ mod.registers.r4\[6\] _0508_ _3237_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_131_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _2924_ _2925_ _2926_ _2917_ _2923_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_77_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _2033_ _2868_ _2875_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3965__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4146__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5646__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4621__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout153_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3890_ _0813_ _0814_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6251__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _2431_ _2432_ _2434_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4511_ _1351_ _1336_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5491_ _2276_ _2379_ _2381_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4137__A1 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _0627_ _1410_ _1411_ _1333_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4137__B2 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4373_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _2802_ _1885_ mod.pc\[7\] _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3324_ _3175_ _3176_ _3163_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6429__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5637__A1 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _2730_ _2069_ _2755_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _0043_ net175 mod.ldr_hzd\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _0377_ net176 mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3820__B1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ mod.registers.r11\[7\] _2607_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6365__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6872__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ mod.registers.r9\[14\] _2562_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _1442_ _1254_ _1513_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5689_ _2422_ _2515_ _2518_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4679__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4300__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__B1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5800__A1 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__C2 _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__B1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6071__I _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6600__I0 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4390__I1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6745__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_340 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_351 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_362 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_373 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6044__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4991_ _1915_ _1950_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6730_ _0234_ net40 mod.registers.r8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6895__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3942_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3802__B1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6661_ _0165_ net92 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3873_ mod.pc_2\[8\] _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5612_ mod.registers.r6\[14\] _2466_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6592_ net3 mod.des.des_dout\[31\] _3142_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5543_ _2253_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3581__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5474_ mod.registers.r4\[6\] _2368_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _0992_ _1394_ _1391_ _1379_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3869__B1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4356_ _1307_ _1314_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3307_ _3158_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4287_ _0551_ _1022_ _1026_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5086__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4833__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6156__I _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6928_ _0026_ net162 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout44 net51 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout55 net63 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6859_ _0360_ net183 mod.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout66 net68 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout77 net79 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout88 net91 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout99 net102 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6618__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4521__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6274__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A2 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4037__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A3 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6015__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3563__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__B2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _1177_ _1179_ _0826_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4512__B2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1861_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ mod.registers.r12\[9\] _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _1038_ _1039_ _1040_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_83_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__A2 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__B1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _1915_ _1933_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ _0217_ net40 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3925_ _0890_ _0892_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6644_ _0148_ net137 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _3133_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3787_ _0728_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4200__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3554__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6910__CLK net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5457_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4408_ _0987_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5388_ _2301_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout201 net202 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout212 net218 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4339_ _0454_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5059__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6009_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3490__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A3 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__I _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6550__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3793__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _0669_ _0528_ _0674_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4981__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _1339_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6933__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3641_ _0609_ _3213_ _3214_ _3218_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_127_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ mod.pc_1\[0\] _2995_ _2996_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3572_ _0448_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ mod.des.des_dout\[30\] _2248_ _2250_ _2252_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ mod.valid1 _2709_ _2151_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5289__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _2169_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _2092_ _2122_ _2129_ _1896_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6238__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4124_ _1076_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4055_ _3226_ _0618_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__B _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6434__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ mod.pc\[1\] _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _0799_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4972__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6627_ _0131_ net138 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3839_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _3118_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ mod.registers.r5\[1\] _2391_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6489_ _3082_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4129__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6806__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__C1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3968__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4191__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5423__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout183_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5860_ _2536_ _2627_ _2632_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _0942_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _2554_ _2585_ _2588_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _1346_ _1335_ _1400_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4673_ _1072_ _1549_ _1642_ _1060_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6203__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6412_ _2141_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3624_ _0576_ _0592_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4706__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _2950_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3555_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6459__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6459__B2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6274_ _2936_ _2937_ _2938_ _2929_ _2935_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3486_ _3234_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4658__B _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ mod.des.des_dout\[21\] _2167_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6829__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _2092_ _2108_ _2113_ _1924_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3693__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3693__B2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4107_ mod.funct3\[0\] _1023_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _2041_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4038_ _1005_ _1006_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6979__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _2712_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6113__B _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__I _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__A1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3920__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5122__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3684__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3684__B2 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4750__C _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__C1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A1 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3340_ mod.instr_2\[17\] _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3911__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5113__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _1971_ _1972_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3675__A1 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6961_ _0059_ net213 mod.des.des_dout\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3427__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__B _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5912_ mod.registers.r13\[6\] _2662_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3978__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3401__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _0393_ net145 mod.instr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ mod.registers.r11\[13\] _2619_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ mod.registers.r10\[3\] _2574_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4725_ _0922_ _1408_ _1693_ _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5328__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4232__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4656_ _1495_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3607_ _3265_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4155__A2 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__A1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ _1401_ _0912_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3902__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3538_ _0418_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6326_ _2955_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ mod.des.des_dout\[11\] _2921_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3469_ _3284_ _0416_ _0425_ _0426_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5208_ _1850_ _2143_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7007__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6188_ mod.pc_1\[7\] _2869_ _2873_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _2095_ _2097_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4407__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3969__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4394__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5591__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5343__A1 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3981__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4298__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5646__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout146_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4385__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5582__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _0776_ _0803_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ mod.registers.r4\[12\] _2380_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4441_ _0790_ _0775_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4137__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3891__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4372_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3896__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _2017_ _2780_ _2812_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3323_ mod.instr_2\[14\] _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _2729_ mod.pc0\[9\] _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5637__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__I0 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3840__B _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout59_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _0042_ net174 mod.ldr_hzd\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4073__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3820__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ _0376_ net192 mod.pc_1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__B2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ _2546_ _2606_ _2610_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _2289_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _1675_ _1676_ _1440_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5688_ mod.registers.r8\[9\] _2516_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4128__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _1468_ _0555_ _1608_ _0623_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5876__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ mod.instr_2\[3\] _2958_ _2963_ mod.instr\[3\] _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4300__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4064__A1 mod.registers.r11\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__B2 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3811__B2 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6697__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6600__I1 mod.des.des_dout\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5316__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_330 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_341 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_352 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_363 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_374 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4990_ _1952_ _1955_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _0908_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3802__B2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6660_ _0164_ net144 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3872_ _0812_ _0827_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5611_ _2436_ _2465_ _2468_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6591_ _3143_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3566__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4763__C1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5542_ _2417_ _2418_ _2420_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5307__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _2218_ _2367_ _2370_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5606__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__B1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4424_ _1376_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5858__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3869__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__B2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ _1315_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3306_ mod.instr_2\[14\] _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ mod.pc_2\[6\] _1205_ _0510_ _0523_ _1047_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_98_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4294__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5794__A1 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _0025_ net182 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3796__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6172__I _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout45 net51 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6858_ _0359_ net191 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout56 net63 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout67 net68 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout78 net79 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5546__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5809_ _2597_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6594__I0 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _0293_ net71 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5516__I _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4521__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3324__A3 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6274__A2 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__A3 _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4037__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__B2 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6585__I0 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4760__A2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4330__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6712__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4140_ _0888_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6265__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4071_ mod.registers.r12\[6\] _0887_ _3211_ mod.registers.r13\[6\] _1041_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6862__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4028__A1 mod.registers.r15\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__B2 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _1916_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6712_ _0216_ net53 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3924_ mod.registers.r2\[4\] _0893_ _3174_ mod.registers.r4\[4\] mod.registers.r10\[4\]
+ _0602_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _0147_ net136 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5528__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6576__I0 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3855_ mod.pc_2\[11\] _0777_ _0819_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3786_ _0683_ _0684_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4200__A1 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ mod.des.des_dout\[24\] net9 _3129_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4200__B2 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _2217_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5456_ _2358_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4407_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5700__A1 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _2236_ _2309_ _2314_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout202 net203 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout213 net215 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4338_ _0683_ _0684_ _0680_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6167__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4269_ _0988_ _0990_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__A3 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6008_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3490__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5020__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4415__I _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6735__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4742__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3702__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3481__A2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ mod.registers.r15\[2\] _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6183__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3571_ _0446_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5930__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5310_ _2213_ _2251_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6290_ _2948_ _2889_ _2949_ _2891_ _2742_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _2136_ _1604_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5172_ _2126_ _2127_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6238__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4123_ _3238_ _1078_ _1088_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4054_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout41_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4235__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4956_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3907_ _0811_ _0842_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_32_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _1849_ mod.instr_2\[3\] _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6626_ _0130_ net140 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6174__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3838_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4185__B1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _3123_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4724__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3769_ mod.registers.r4\[12\] _0738_ _3266_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6488_ mod.des.des_dout\[5\] net3 _3080_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _2261_ _2343_ _2347_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4488__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3314__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5988__A1 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3999__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__C2 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5912__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4191__A3 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout176_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6900__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4810_ _1390_ _1778_ _1779_ _1392_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5790_ mod.registers.r10\[9\] _2586_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _1328_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4672_ _1072_ _0944_ _0938_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6411_ _1849_ _2883_ _3028_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3623_ _0495_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4706__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5903__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3509__A3 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6342_ _2707_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3554_ mod.pc_2\[6\] _0499_ _0510_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6273_ mod.des.des_dout\[15\] _2933_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3485_ _3254_ _3180_ _3222_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _3263_ _2168_ _2170_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5131__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout89_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _2092_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3693__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4106_ _0591_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5086_ _1970_ _2040_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4037_ mod.registers.r11\[7\] _0605_ _3199_ mod.registers.r9\[7\] _1007_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _2711_ _1884_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4939_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _0113_ net139 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3309__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6556__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3684__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4881__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6923__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4633__A1 _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4149__B1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__C2 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A3 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3675__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3889__I _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _0058_ net216 mod.des.des_dout\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3427__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ _2407_ _2661_ _2664_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _0392_ net147 mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ _2560_ _2618_ _2620_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5773_ _2536_ _2572_ _2577_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4724_ _0526_ _1103_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4655_ _1260_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3606_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A2 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4586_ _1555_ _0454_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6325_ _2971_ _2974_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3537_ mod.registers.r11\[6\] _0505_ _0506_ mod.registers.r2\[6\] _0507_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _2718_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A2 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3468_ mod.registers.r15\[0\] _0435_ _0437_ mod.registers.r12\[0\] _0438_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6946__CLK net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ mod.rd_3\[0\] _2144_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6187_ _2017_ _2868_ _2874_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3399_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A1 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _0957_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5069_ _1911_ _2004_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4615__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3969__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3748__B _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5591__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A3 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5203__B _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4606__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4909__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout139_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _1409_ _0827_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6531__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3345__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ _0621_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3896__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6110_ _2767_ _2811_ _2778_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ mod.instr_2\[15\] _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__I1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3412__I _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _0041_ net166 mod.ldr_hzd\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4073__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6874_ _0375_ net185 mod.pc_1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3820__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3568__B _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5825_ mod.registers.r11\[6\] _2607_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5756_ _2564_ _2561_ _2565_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _1515_ _1252_ _1249_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ _2417_ _2515_ _2517_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _1316_ _0576_ _0592_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6522__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4569_ _1538_ _0724_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5089__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ mod.instr\[7\] _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__A1 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3322__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4064__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3811__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5564__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3992__I _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5712__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_320 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_331 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_342 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_353 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_364 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_375 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3940_ _3227_ _0902_ _0909_ _0903_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_32_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3802__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _0828_ _0553_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5610_ mod.registers.r6\[13\] _2466_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6590_ net2 mod.des.des_dout\[30\] _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3566__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4763__B1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5541_ mod.registers.r5\[8\] _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3566__B2 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__C2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5472_ mod.registers.r4\[5\] _2368_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5307__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3318__A1 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4423_ _1391_ _1380_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3318__B2 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3869__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4354_ _1317_ _1319_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3305_ mod.instr_2\[15\] _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4285_ _1249_ _1252_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6024_ _2706_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout71_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A1 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5243__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4046__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _0024_ net163 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _0358_ net182 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout46 net47 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout57 net62 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout68 net74 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5808_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout79 net82 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6788_ _0292_ net135 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4349__A3 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6594__I1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5739_ _2550_ _2551_ _2553_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6402__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3317__I _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4285__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5482__A1 mod.registers.r4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5707__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3720__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6538__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ mod.registers.r14\[6\] _3208_ _3169_ mod.registers.r7\[6\] _1040_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5473__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__A2 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A1 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4972_ _1051_ _1935_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _0215_ net53 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5110__C _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3923_ _3191_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6642_ _0146_ net136 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3854_ _0820_ _0821_ _0822_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5528__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6576__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3539__A1 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _3132_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3785_ _0727_ _0728_ _0740_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5617__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4200__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _2403_ _2404_ _2406_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5455_ _2356_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4406_ _1245_ _1247_ _1303_ _1304_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5386_ mod.registers.r2\[7\] _2310_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5700__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout203 mod.clk net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4337_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6687__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4268_ _1225_ _1230_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5464__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6007_ _2711_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4806__A4 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4199_ mod.registers.r11\[11\] _0705_ _0697_ mod.registers.r1\[11\] _1169_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _0007_ net142 mod.instr_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3702__B2 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3510__I _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6042__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout121_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout219_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3570_ mod.registers.r15\[7\] _0435_ _0437_ mod.registers.r12\[7\] _0540_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5930__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _2182_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _2126_ _2127_ _2056_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _0615_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A1 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4249__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4053_ _3232_ _3251_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_in[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3420__I _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _1895_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _0802_ _0860_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ mod.instr_2\[4\] mod.instr_2\[3\] _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6625_ _0129_ net139 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3837_ _0804_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6174__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4185__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ mod.des.des_dout\[16\] net19 _3119_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3768_ _0419_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5921__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _2185_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _3081_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3699_ mod.pc_2\[1\] _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5438_ mod.registers.r3\[10\] _2344_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4488__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6178__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5369_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5810__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__B2 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4176__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3518__A4 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5428__A1 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4100__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6037__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout169_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__A1 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _1352_ _1630_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__B1 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ _1315_ _1314_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4167__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ mod.rd_3\[1\] _2884_ _3017_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3622_ _0579_ _0591_ _3262_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _2978_ _2984_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3553_ _0513_ _0516_ _0519_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _2718_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3484_ _3246_ _3262_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5667__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ mod.pc_2\[12\] _1089_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_69_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5419__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4105_ _0578_ _1074_ _0896_ _0898_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__3693__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5085_ _1970_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5630__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6092__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4036_ mod.registers.r2\[7\] _0701_ _3195_ mod.registers.r10\[7\] _1006_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6725__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ net12 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6395__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6461__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6875__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4938_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _1814_ _1835_ _1015_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6608_ _0112_ net130 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3905__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6539_ _3094_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5658__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4881__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5540__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4584__C _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4633__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6572__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__B2 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5715__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__C1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__B2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6748__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5821__A1 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ mod.registers.r13\[5\] _2662_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6890_ _0391_ net145 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5841_ mod.registers.r11\[12\] _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4388__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ mod.registers.r10\[2\] _2574_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _1675_ _1669_ _1484_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _1071_ _1267_ _1056_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5888__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3605_ _0556_ _0557_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4585_ _1265_ _1070_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6324_ _1391_ _2968_ _2972_ mod.instr\[8\] _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4560__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3536_ _0411_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6255_ mod.instr\[11\] _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3467_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4312__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _1849_ _2143_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6186_ mod.pc_1\[6\] _2869_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3398_ _3230_ _3231_ mod.instr_2\[1\] _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5137_ mod.funct7\[0\] _1206_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5360__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6065__A1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _2005_ _2024_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4019_ _0799_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3823__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A1 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3339__C1 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6540__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4146__A4 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6366__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A3 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A3 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__A2 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6531__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout201_I net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ _3173_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6477__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _2752_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__C1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6942_ _0040_ net165 mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4073__A3 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6873_ _0374_ net185 mod.pc_1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _2544_ _2606_ _2609_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5755_ mod.registers.r9\[13\] _2562_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3584__A2 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _0526_ _1103_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5686_ mod.registers.r8\[8\] _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6913__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4637_ _1572_ _1605_ _1606_ _1515_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4568_ _0899_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6307_ _2950_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3519_ _3252_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1468_ _1305_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A1 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _2908_ _2901_ _2910_ _2905_ _2911_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4836__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _1893_ _2859_ _2862_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6119__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4049__B1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__A2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3732__C1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A2 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_310 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_321 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6029__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_332 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_343 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_354 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_365 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_376 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout151_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3870_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6936__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _2390_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3566__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__B2 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _2205_ _2367_ _2369_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4422_ _0914_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3318__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4353_ _1317_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3304_ _3157_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4284_ _1253_ _1093_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _2739_ _2740_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3423__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout64_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4963__B _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__A3 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ _0023_ net163 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _0357_ net189 mod.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout47 net50 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout58 net62 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5807_ _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4203__B1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout69 net73 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6787_ _0291_ net124 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3999_ mod.registers.r6\[15\] _0966_ _0967_ mod.registers.r5\[15\] _0968_ mod.registers.r8\[15\]
+ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5738_ mod.registers.r9\[8\] _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _2394_ _2502_ _2506_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4506__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3333__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3493__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6791__D _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5234__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6431__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3489__B _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__B1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3508__I _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout199_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3484__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5225__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4971_ _1917_ _1937_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6710_ _0214_ net59 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3922_ mod.registers.r14\[4\] _0891_ _0705_ mod.registers.r11\[4\] _0892_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3853_ mod.registers.r13\[11\] _0520_ _0521_ mod.registers.r1\[11\] _0823_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6641_ _0145_ net136 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4736__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3539__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _0742_ _0744_ _0750_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6572_ mod.des.des_dout\[23\] net8 _3129_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5523_ mod.registers.r5\[4\] _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5454_ _2155_ _2157_ _2159_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4405_ _1326_ _1330_ _1348_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3862__B _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5161__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _2229_ _2309_ _2313_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4336_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout204 net205 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout215 net217 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4267_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6006_ _2724_ _2727_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5464__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4198_ mod.registers.r14\[11\] _0891_ _0703_ mod.registers.r9\[11\] mod.registers.r2\[11\]
+ _0893_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_83_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6908_ _0409_ net142 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _0340_ net156 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5152__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6631__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3702__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3466__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3998__I _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5718__I _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4194__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout114_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__I _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5170_ mod.pc_2\[13\] _0955_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4121_ _1089_ _1090_ _0617_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5446__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _3254_ _1008_ _1020_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_96_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3457__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput4 io_in[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4957__A1 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _1900_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3905_ _0828_ _0861_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_32_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4885_ mod.ldr_hzd\[3\] _1852_ _1854_ mod.ldr_hzd\[1\] _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _0128_ net93 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3836_ _0577_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4185__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _3122_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3767_ mod.registers.r11\[12\] _0735_ _0736_ mod.registers.r2\[12\] _0737_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6654__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5506_ _2386_ _2389_ _2392_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6486_ mod.des.des_dout\[4\] net2 _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3698_ _0650_ _0666_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5134__A1 mod.pc_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5437_ _2254_ _2343_ _2346_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5368_ _2300_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3696__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4319_ _0731_ _0734_ _0737_ _0739_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5299_ _1951_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3999__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5538__I _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5373__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3687__A1 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4100__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5600__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _1420_ _1632_ _1634_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _0580_ _0421_ _0585_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4167__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ mod.registers.r13\[6\] _0520_ _0521_ mod.registers.r1\[6\] _0522_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6340_ _1136_ _2982_ _2979_ mod.instr\[14\] _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6271_ mod.instr\[15\] _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5116__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3483_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _2171_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3678__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4875__B1 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4875__C2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5153_ _2094_ _2098_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4104_ _0567_ _0572_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _0843_ _2042_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_96_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6092__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4035_ mod.registers.r15\[7\] _0963_ _3186_ mod.registers.r6\[7\] _3189_ mod.registers.r5\[7\]
+ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_65_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3431__I mod.instr_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ mod.valid0 _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ mod.des.des_counter\[0\] _3150_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _1833_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5355__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6607_ _0111_ net130 mod.registers.r1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3819_ _0784_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4799_ _1665_ _1360_ _1367_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6538_ _3092_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__B1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _1819_ _3064_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3606__I _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3669__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5594__A1 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__B1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__C2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4321__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__I _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A3 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _2600_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4388__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5585__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5771_ _2534_ _2572_ _2576_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3596__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4722_ _1675_ _1670_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4653_ _1445_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5906__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3604_ _0567_ _0572_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4584_ _1517_ _1522_ _1523_ _1553_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3899__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3899__B2 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6323_ _2971_ _2973_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3535_ _3290_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3426__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _2920_ _2913_ _2922_ _2917_ _2923_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3466_ _3281_ _0417_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ mod.rd_3\[1\] _2144_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4312__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3397_ _3244_ _3247_ _3249_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6185_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5136_ mod.pc_2\[11\] _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _1790_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6842__CLK net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _0950_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3823__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3823__B2 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6992__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A2 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2680_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3339__B1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3339__C2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__I0 mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3354__A3 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3336__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4303__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5551__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6056__A2 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6583__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4909__A4 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5319__A1 mod.des.des_dout\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5726__I _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6715__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3345__A3 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3320_ _3166_ _3168_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_125_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3502__B1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3502__C2 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _0039_ net197 mod.ldr_hzd\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3805__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6292__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _0373_ net192 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5823_ mod.registers.r11\[5\] _2607_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5754_ _2283_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4705_ _0526_ _1103_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4781__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5685_ _2503_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _1454_ _1448_ _1453_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5730__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _1401_ _0623_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6306_ _2759_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3518_ _0472_ _0474_ _0475_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_103_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _0691_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6237_ _2788_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3449_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ mod.pc_1\[0\] _2861_ _2822_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _2060_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4049__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6099_ _1389_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4049__B2 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5549__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A3 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6210__A2 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6888__CLK net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__B1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__C2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__I _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4288__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_300 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_311 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_322 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_333 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_344 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_355 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_366 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3799__B1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout144_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3685__B _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3971__B1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5470_ mod.registers.r4\[4\] _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ _3229_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4352_ _1320_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3303_ mod.des.des_counter\[2\] _3151_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4283_ _0591_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ _2726_ _1983_ _2731_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout57_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _0022_ net164 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ _0356_ net158 mod.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout48 net50 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _2327_ _2499_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout59 net62 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4203__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _0290_ net134 mod.registers.r12\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3998_ _0473_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4203__B2 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5737_ _2531_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5951__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5668_ mod.registers.r8\[1\] _2504_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5703__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _0938_ _1588_ _1061_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5599_ _2417_ _2459_ _2461_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6503__I0 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__B2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6195__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5276__I _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5942__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5170__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5225__B _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1206_ _0492_ _1045_ _0669_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__4433__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ _3208_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _0144_ net92 mod.registers.r3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3852_ mod.registers.r5\[11\] _0517_ _0518_ mod.registers.r7\[11\] _0822_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5933__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _3131_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3783_ mod.registers.r9\[12\] _0751_ _0752_ mod.registers.r3\[12\] _0753_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5186__I _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5522_ _2390_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _2355_ _2149_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4404_ _0992_ _1349_ _1361_ _1368_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5384_ mod.registers.r2\[6\] _2310_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5161__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4335_ _0808_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout205 net207 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3434__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout216 net217 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4266_ _1004_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _2726_ _1903_ _0003_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _1165_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _0408_ net168 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6838_ _0339_ net161 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4188__B1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4727__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5924__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _0273_ net134 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5152__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3344__I mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6101__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3466__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6404__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A1 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3519__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__B2 mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ mod.funct7\[1\] _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4051_ _3264_ _1002_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4654__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 io_in[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__B2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _1890_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4884_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _0127_ net93 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3835_ _0560_ _0618_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ mod.des.des_dout\[15\] net18 _3119_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3766_ _0412_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ mod.registers.r5\[0\] _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ _3074_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3697_ _0528_ _0552_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_118_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ mod.registers.r3\[9\] _2344_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5134__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5367_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3696__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4318_ _1226_ _1202_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5298_ _2208_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ _1152_ _1218_ _1143_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4645__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5819__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3687__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6086__B1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6389__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5729__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A2 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3620_ _0586_ _0587_ _0588_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4167__A3 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3551_ _0448_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _2932_ _2925_ _2934_ _2929_ _2935_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5116__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3482_ _3263_ _3266_ _0423_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4175__I0 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5221_ _1792_ _3257_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4875__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4875__B2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5152_ mod.pc_2\[11\] _2097_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4103_ _1056_ _1060_ _1064_ _1071_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _2043_ _2028_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4627__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _0779_ _1003_ _0789_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3850__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5985_ _1895_ _1884_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5639__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6621__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4936_ _3224_ _1905_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4867_ _1820_ _1834_ _1835_ _1819_ _1836_ _1818_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_6606_ _0110_ net129 mod.registers.r1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3818_ _0785_ _0786_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5355__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _1352_ _1324_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6537_ _2427_ _3106_ _3111_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3905__A3 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3749_ _0595_ _0699_ _0710_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_4_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6304__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _3068_ _3069_ _3057_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6304__B2 mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5419_ _2194_ _2330_ _2335_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ net20 _2152_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3669__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4094__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__B _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6543__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3357__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5284__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4857__B2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3532__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A4 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout174_I net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6644__CLK net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6064__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ mod.registers.r10\[1\] _2574_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3596__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6794__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4721_ _1689_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3596__B2 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _1580_ _1261_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6534__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3348__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3603_ mod.pc_2\[4\] _0499_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4312__B _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4583_ _1331_ _1543_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _1392_ _2968_ _2972_ mod.instr\[7\] _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3534_ mod.registers.r14\[6\] _0502_ _0503_ mod.registers.r6\[6\] _0504_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4560__A3 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _2741_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3465_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5204_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout87_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6184_ _2752_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _3248_ _3228_ mod.funct3\[0\] _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_97_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ _2093_ _2080_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3442__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ mod.pc_2\[7\] _2025_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__B _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__A1 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _3247_ _0958_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3823__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5369__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5968_ _2427_ _2694_ _2699_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4379__A3 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4919_ _1885_ _1887_ mod.valid0 _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5899_ _2385_ _2654_ _2657_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6525__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3339__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3339__B2 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6128__I1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5500__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3511__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__A1 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5567__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__C1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3593__A4 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4358__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3502__A1 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3502__B2 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _0038_ net195 mod.rd_3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _0372_ net185 mod.pc_1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5007__A1 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5822_ _2540_ _2606_ _2608_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3569__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5753_ _2560_ _2561_ _2563_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5917__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4230__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _1654_ _1657_ _1658_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _2501_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _1300_ _0940_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1501_ _1419_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_116_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _2760_ _2960_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _0479_ _0481_ _0484_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4497_ _0726_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6236_ mod.des.des_dout\[6\] _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3448_ _0415_ _0416_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_131_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4297__A2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _3230_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _2059_ _2061_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6098_ _2783_ _2791_ _2798_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4049__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5049_ _2008_ _2009_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5549__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3980__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__B1 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3732__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3732__B2 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5562__I _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4288__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5485__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A4 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6594__S _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_301 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_312 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_323 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_334 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_345 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_356 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_367 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3799__B2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4212__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5737__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout137_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3971__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3971__B2 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _3227_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3723__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _0579_ _0525_ _0681_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3302_ _3156_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4282_ _1250_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6982__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _2723_ mod.pc0\[4\] _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _0021_ net163 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6854_ _0355_ net158 mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _2568_ _2591_ _2596_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6785_ _0289_ net134 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5400__A1 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _0468_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4203__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _2529_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _2386_ _2502_ _2505_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _1056_ _1549_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5703__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ mod.registers.r6\[8\] _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4549_ _1518_ _1514_ _1075_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6503__I1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5467__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6219_ mod.des.des_dout\[2\] _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3786__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5557__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6855__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3705__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3705__B2 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5292__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3484__A3 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__B _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ mod.registers.r12\[4\] _0888_ _0889_ mod.registers.r13\[4\] _0890_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3851_ mod.registers.r9\[11\] _0511_ _0512_ mod.registers.r3\[11\] _0821_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4371__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4197__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6570_ mod.des.des_dout\[22\] net7 _3129_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3782_ _0512_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5933__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _2388_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6499__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _2146_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5697__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _0990_ _1369_ _1372_ _1246_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6298__I _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5383_ _2218_ _2309_ _2312_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4334_ _1298_ _1299_ _3241_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout206 net207 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout217 net218 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6497__I0 mod.des.des_dout\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4265_ _3247_ _1231_ _1232_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6004_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4196_ _1161_ _1164_ _0839_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_39_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3450__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _0407_ net168 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4975__A3 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _0338_ net156 mod.pc0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4281__I _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4188__B2 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5924__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6768_ _0272_ net112 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5719_ mod.registers.r9\[3\] _2532_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6699_ _0203_ net39 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A1 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3625__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__I _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4360__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5840__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5860__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3360__I _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3535__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4351__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4103__B2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ _1009_ _1018_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_37_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4654__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ mod.pc0\[1\] _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3903_ _0862_ _0464_ _0867_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6159__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ mod.instr_2\[4\] _1850_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3834_ _3253_ _0599_ _0613_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_60_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _0126_ net131 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3917__A1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _3121_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3765_ _3291_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__C _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6484_ _3079_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3696_ _0651_ _0464_ _0656_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _2245_ _2343_ _2345_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5366_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4893__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4317_ _1276_ _1286_ _1223_ _1203_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_102_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5297_ _2191_ _2040_ _2209_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4248_ _1213_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5842__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3448__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4276__I _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4179_ _0858_ _1147_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3853__B1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3355__I _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5570__I _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6086__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__B1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__A1 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6389__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4167__A4 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout217_I net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3550_ _0446_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3481_ _0432_ _0438_ _0443_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5220_ mod.ins_ldr_3 mod.valid_out3 net15 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4175__I1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4875__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _1987_ _2108_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4102_ _1062_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5082_ _0530_ _2025_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4627__A2 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _0687_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_84_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2708_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _3225_ _1387_ _1903_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4866_ _1135_ _1136_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__CLK net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6605_ _0109_ net129 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3817_ mod.registers.r14\[14\] _0732_ _0730_ mod.registers.r10\[14\] _0787_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4012__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _1345_ _1481_ _1638_ _1467_ _1660_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3748_ _0624_ _0693_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6536_ mod.registers.r15\[11\] _3107_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _3055_ _3036_ _3066_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3679_ _0644_ _0645_ _0646_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6304__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ mod.registers.r3\[2\] _2332_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6398_ _2152_ _3020_ _2831_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3669__A3 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5349_ _2168_ _2136_ _1435_ _2273_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4618__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A1 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5291__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6435__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5565__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4003__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4554__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4609__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__A1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4085__A3 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout167_I net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4720_ _1467_ _1421_ _1540_ _1566_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3596__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _1607_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6534__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3602_ _0568_ _0569_ _0570_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4545__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ _1367_ _1546_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6321_ _2962_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3533_ _3286_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6252_ mod.des.des_dout\[10\] _2921_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ _0429_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5203_ _3244_ _2152_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6183_ _1999_ _2868_ _2871_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3395_ _3226_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5134_ mod.pc_2\[10\] _0958_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _2026_ _2012_ _2027_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _0687_ _0984_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ mod.registers.r14\[11\] _2695_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4918_ net13 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4784__B2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ mod.registers.r13\[0\] _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4849_ mod.ldr_hzd\[14\] _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3339__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _3094_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4729__I _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3633__I _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3511__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6213__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__C2 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5295__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3808__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3971__C _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3502__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6452__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6761__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3805__A3 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4374__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _0371_ net192 mod.pc_1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ mod.registers.r11\[4\] _2607_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3569__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ mod.registers.r9\[12\] _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4230__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ _1664_ _1668_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _2414_ _2509_ _2514_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4518__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4634_ _1585_ _1586_ _1590_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4565_ _1532_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5191__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6304_ _0903_ _2958_ _2951_ mod.instr\[2\] _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3516_ mod.registers.r15\[1\] _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4496_ _3242_ _1461_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6235_ _2888_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3447_ _3270_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5494__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3378_ mod.instr_2\[0\] _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6166_ _2856_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _2076_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6097_ _1980_ _2766_ _2800_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6443__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5048_ mod.pc_2\[5\] _1991_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input12_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6999_ _0097_ net207 mod.des.des_dout\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4757__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3980__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5182__B2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6634__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4459__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3363__I _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5485__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__C1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5999__B _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4532__I1 _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_302 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_313 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_324 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_335 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_346 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_357 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_368 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3799__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3538__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3971__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4797__C _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4350_ _0757_ _0861_ _0551_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3723__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3301_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _0574_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _2708_ _2738_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6425__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ _0020_ net164 mod.pc_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__A3 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _0354_ net159 mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5804_ mod.registers.r10\[15\] _2592_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout39 net42 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_6784_ _0288_ net113 mod.registers.r12\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _0600_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5400__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5735_ _2244_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5666_ mod.registers.r8\[0\] _2504_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5164__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4617_ _1306_ _1407_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5663__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ _2447_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _1073_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4479_ _0812_ _1069_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _2888_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4675__B1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6494__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6149_ _2816_ _2837_ _2841_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5219__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6416__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4978__A1 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5059__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3705__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4130__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A1 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3641__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3641__B2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3850_ mod.registers.r15\[11\] _0514_ _0515_ mod.registers.r12\[11\] _0820_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3781_ _0511_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5394__A1 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5146__A1 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _2296_ _2349_ _2354_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__B _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5697__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4402_ _0988_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5382_ mod.registers.r2\[5\] _2310_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4099__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4333_ _1298_ _1299_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5449__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout207 net208 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout218 net219 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4264_ _0926_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _2711_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4195_ _0839_ _1161_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3731__I _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout62_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3880__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _0406_ net173 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _0337_ net154 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5385__A1 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4188__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6767_ _0271_ net115 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3979_ _3243_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4727__A4 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5718_ _2198_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ _0202_ net53 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5649_ _2472_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__I1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5860__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3871__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4472__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__A1 mod.registers.r2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4351__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6479__I1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3551__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout197_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__A1 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4951_ _1915_ _1910_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5478__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3614__A1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3902_ _0868_ _0869_ _0870_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_32_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4315__C _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6621_ _0125_ net131 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3833_ _0790_ _0800_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ mod.des.des_dout\[14\] net17 _3119_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3764_ mod.registers.r14\[12\] _0732_ _0733_ mod.registers.r6\[12\] _0734_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5503_ _2387_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6316__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ mod.des.des_dout\[3\] net19 _3075_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3726__I _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3695_ _0657_ _0658_ _0659_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5434_ mod.registers.r3\[8\] _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4342__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _2150_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4316_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ mod.pc_2\[8\] _2221_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4247_ _1214_ _1215_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3461__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6845__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4178_ _0858_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3853__A1 mod.registers.r13\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3853__B2 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4506__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3605__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5388__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6995__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__B1 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5358__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6819_ _0323_ net123 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4467__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__B2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4636__A3 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7000__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5298__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5349__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__I _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3780__B1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout112_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ mod.registers.r13\[0\] _0447_ _0449_ mod.registers.r1\[0\] _0450_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6868__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _2107_ _1489_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6078__B mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4101_ _1068_ _0929_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5081_ _0530_ _2025_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4032_ mod.funct7\[2\] _0614_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3835__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A1 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ _2708_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5052__A3 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3599__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4934_ _3155_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _0480_ _3256_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6604_ _0108_ _0003_ net206 mod.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3816_ mod.registers.r13\[14\] _0745_ _0738_ mod.registers.r4\[14\] _0733_ mod.registers.r6\[14\]
+ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4012__A1 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1760_ _1761_ _3243_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6535_ _2424_ _3106_ _3110_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3747_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3456__I mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6466_ _1818_ _3064_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3678_ mod.registers.r13\[2\] _0541_ _0542_ mod.registers.r1\[2\] _0647_ _0648_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4315__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _2186_ _2330_ _2334_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6397_ mod.valid_out3 _2153_ _2713_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ _2270_ _2284_ _2285_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3405__B _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _0902_ _0561_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__I _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4251__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4003__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4003__B2 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3357__A3 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3366__I mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4306__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3817__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3817__B2 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6361__B _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _0918_ _1614_ _1615_ _1616_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[18] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3601_ mod.registers.r5\[4\] _0440_ _3292_ mod.registers.r11\[4\] _0571_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4545__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5742__A1 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3348__A3 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _1547_ _1549_ _1550_ _1098_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6690__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _2759_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3532_ _3282_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6251_ _2888_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3463_ _3281_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3505__B1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5202_ net12 _2142_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6182_ mod.pc_1\[5\] _2869_ _2864_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3394_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _2005_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _2008_ _2009_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6470__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _0955_ _0561_ _0720_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4481__A1 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4233__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5966_ _2424_ _2694_ _2698_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4917_ _1886_ _1883_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4784__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2655_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4848_ mod.ldr_hzd\[13\] _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5733__A1 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _1165_ _1485_ _1369_ _1185_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ _3092_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _2715_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3914__I _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3511__A3 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__B2 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5724__A1 mod.registers.r9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4160__B1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6906__CLK net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__S _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _2600_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _2531_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3569__A3 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4702_ _1128_ _1669_ _1573_ _1330_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5682_ mod.registers.r8\[7\] _2510_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4633_ _1596_ _1601_ _1602_ _0917_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4518__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _1362_ _1533_ _0812_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6303_ _2760_ _2959_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3515_ _3181_ _3197_ _3158_ _3184_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_104_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4495_ _1302_ _1464_ _1246_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6234_ mod.instr\[6\] _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3446_ _3285_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3377_ mod.instr_2\[2\] _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _2075_ _0958_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _2767_ _2799_ _2778_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _2010_ _1994_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4454__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ _0096_ net214 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5954__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5949_ _2680_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3909__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6929__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__C2 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4693__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_303 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_314 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_325 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_336 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_347 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_358 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_369 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5945__A1 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3708__B1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5173__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3300_ _3153_ _3154_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4280_ _3245_ _0896_ _0898_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_113_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _0019_ net168 mod.pc_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _0353_ net157 mod.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6189__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5803_ _2566_ _2591_ _2595_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4334__B _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4739__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ _0287_ net116 mod.registers.r12\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5936__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ mod.registers.r12\[15\] _0962_ _0964_ mod.registers.r15\[15\] _0965_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _2548_ _2541_ _2549_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _1572_ _1582_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5164__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6361__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _2445_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _1513_ _1516_ _1301_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4478_ _1445_ _1446_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6217_ mod.instr\[2\] _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ _3275_ _3277_ _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4675__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3478__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__B2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _2102_ _2824_ _2844_ _2789_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6416__A2 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6079_ _1943_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3650__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5854__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6751__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3374__I _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6104__A1 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4115__B1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4969__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A1 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout142_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ mod.registers.r13\[12\] _0745_ _0746_ mod.registers.r1\[12\] _0749_ _0750_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_20_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ mod.registers.r3\[15\] _2350_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4401_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5381_ _2205_ _2309_ _2311_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4332_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout208 net209 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout219 net1 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4263_ _1113_ _0953_ _0957_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_99_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _2723_ mod.pc0\[0\] _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _3245_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5004__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4843__I mod.ldr_hzd\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _0405_ net177 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ _0336_ net153 mod.pc0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6766_ _0270_ net115 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3978_ _3250_ _0463_ _0919_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ _2536_ _2530_ _2537_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6697_ _0201_ net40 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5674__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5648_ _2428_ _2486_ _2491_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5137__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5579_ _2386_ _2446_ _2449_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3320__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__A1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3926__A3 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A3 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4639__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3311__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 io_in[16] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4950_ _1916_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3614__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3901_ mod.registers.r5\[9\] _0547_ _0548_ mod.registers.r7\[9\] _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6797__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6620_ _0124_ net84 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3832_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4024__C1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _3120_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3763_ _0503_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5502_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6482_ _3078_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6316__A1 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3694_ mod.registers.r13\[3\] _0541_ _0542_ mod.registers.r1\[3\] _0663_ _0664_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5433_ _2331_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5364_ _2159_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _1182_ _1278_ _1282_ _1274_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4838__I _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5295_ _2163_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6258__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4246_ mod.registers.r8\[12\] _0968_ _0981_ mod.registers.r9\[12\] _1216_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _1144_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3853__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3605__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6818_ _0322_ net120 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _0253_ net111 mod.registers.r10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__A1 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3652__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4097__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4416__C _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3780__A1 mod.registers.r13\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3780__B2 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout105_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3562__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4100_ _0688_ _0689_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5080_ _1135_ _0954_ _0957_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5285__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ mod.registers.r12\[14\] _0962_ _0996_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_84_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3835__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5037__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _2708_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3599__A1 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1797_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3599__B2 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6537__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _3160_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3815_ mod.registers.r11\[14\] _0735_ _0746_ mod.registers.r1\[14\] _0785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6603_ _3149_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _1699_ _1764_ _1247_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4012__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ mod.registers.r15\[10\] _3107_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _3065_ _3067_ _3057_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3677_ _0609_ _0433_ _0417_ _0563_ _0610_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6812__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ mod.registers.r3\[1\] _2332_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _0758_ _2953_ _3019_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4568__I _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3523__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ mod.registers.r1\[13\] _2277_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3472__I _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6068__A3 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ _2008_ _2210_ _2208_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ _1197_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5399__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4251__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4003__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3514__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3817__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__C1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3557__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6835__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3600_ mod.registers.r12\[4\] _0437_ _0428_ mod.registers.r9\[4\] _0570_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput11 io_in[1] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _1547_ _0944_ _0938_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5742__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3531_ mod.registers.r8\[6\] _3272_ _0500_ mod.registers.r10\[6\] _0501_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6250_ mod.instr\[10\] _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3462_ mod.registers.r9\[0\] _0428_ _0431_ mod.registers.r3\[0\] _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6985__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3505__A1 mod.registers.r11\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5201_ _1886_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4702__B1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6181_ _1980_ _2868_ _2870_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3393_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5132_ _2056_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__B1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ mod.pc_2\[6\] _2009_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _0970_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4481__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ mod.registers.r14\[10\] _2695_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5430__A1 mod.registers.r3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ mod.valid2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5896_ _2652_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4847_ mod.ldr_hzd\[12\] _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4778_ _1384_ _1740_ _1742_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ _0695_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6517_ _2399_ _3093_ _3099_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _3055_ _3044_ _3037_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5497__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6379_ _2713_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5249__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3511__A4 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4224__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__CLK net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3377__I mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4527__A3 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__B1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__B1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4001__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4160__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__B2 mod.registers.r13\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A3 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout172_I net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5767__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4846__S0 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ _2529_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5963__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4701_ _1126_ _1371_ _1670_ _1186_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5681_ _2411_ _2509_ _2513_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4632_ _0901_ _1564_ _1566_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ _0828_ _0553_ _0773_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3514_ _0482_ _0483_ mod.registers.r13\[1\] _0477_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6302_ _1792_ _2958_ _2951_ mod.instr\[1\] _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4494_ _1224_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6233_ _2906_ _2901_ _2907_ _2905_ _2898_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3445_ _3284_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _2857_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout85_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3376_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ mod.pc_2\[10\] _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _2792_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3750__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ mod.pc_2\[5\] _1991_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5651__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _0095_ net209 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _2399_ _2681_ _2687_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5879_ mod.registers.r12\[10\] _2641_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A3 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6301__I _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4142__A1 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__B2 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5890__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_304 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_315 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_326 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_337 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_348 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_359 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6211__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5633__A1 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _0018_ net163 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _0352_ net157 mod.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6189__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5802_ mod.registers.r10\[14\] _2592_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6782_ _0286_ net115 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5936__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3947__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ mod.registers.r9\[7\] _2542_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _2500_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4615_ _1300_ _1582_ _1584_ _3250_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4350__B _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5595_ _2414_ _2453_ _2458_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6361__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4546_ _1249_ _1515_ _1252_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4477_ _0716_ _1310_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5960__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6216_ _2893_ _2719_ _2894_ _2892_ _2855_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3428_ mod.instr_2\[13\] _3268_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5872__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _2842_ _2843_ _2818_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3359_ mod.registers.r12\[0\] _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3883__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6078_ _2768_ _2004_ mod.pc\[2\] _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5624__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5029_ _1992_ _1975_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3650__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3938__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3655__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__B2 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__B _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__B1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5918__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout135_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3565__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ _0932_ _0936_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4354__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ mod.registers.r2\[4\] _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4262_ _0779_ _0789_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout209 net219 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4193_ _0953_ _1091_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3865__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A3 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3617__B1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5082__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ _0404_ net177 mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout48_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__I _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _0335_ net161 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6919__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6765_ _0269_ net111 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3977_ _0922_ _0928_ _0941_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ mod.registers.r9\[2\] _2532_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _0200_ net55 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ mod.registers.r7\[11\] _2487_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ mod.registers.r6\[0\] _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4529_ _1496_ _1497_ _1383_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5845__A1 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__I _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3385__I _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5836__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3698__I0 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__I mod.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3847__B1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3311__A2 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 io_in[17] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_36_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5064__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ mod.registers.r9\[9\] _0544_ _0545_ mod.registers.r3\[9\] _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _3255_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6013__A1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3831_ _0690_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4024__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4024__C2 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ mod.des.des_dout\[13\] net16 _3119_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3762_ _0502_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ mod.des.des_dout\[2\] net18 _3075_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6316__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3693_ _0660_ _0433_ _0661_ _0563_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_9_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4327__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _2329_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6600__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _2154_ _2157_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4314_ _0826_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5294_ _2201_ _2236_ _2237_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5827__A1 mod.registers.r11\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4245_ mod.registers.r6\[12\] _0966_ _0967_ mod.registers.r5\[12\] _1215_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _3266_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__I mod.ldr_hzd\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6741__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _0321_ net121 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5685__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__CLK net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6748_ _0252_ net48 mod.registers.r9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ _0183_ net55 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4318__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4869__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3933__I _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__A2 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4006__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5349__A3 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4557__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4004__I _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4939__I _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6614__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ _0997_ _0998_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3296__A1 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__B _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4245__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5981_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ mod.pc0\[0\] _1892_ _1898_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3599__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4623__B _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _1817_ _1832_ _0478_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6537__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ net8 mod.des.des_dout\[36\] _3136_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3814_ _0780_ _0781_ _0782_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4794_ _1273_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _2421_ _3106_ _3109_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3745_ _3246_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _3055_ _1862_ _3066_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3676_ mod.registers.r9\[2\] _0544_ _0545_ mod.registers.r3\[2\] _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _2177_ _2330_ _2333_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6395_ mod.pc_1\[13\] _2720_ _3017_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3523__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__C _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4720__B2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _2221_ _2007_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4228_ mod.registers.r11\[13\] _0974_ _0972_ mod.registers.r10\[13\] mod.registers.r4\[13\]
+ _0971_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ mod.registers.r12\[8\] _1110_ _0879_ mod.registers.r7\[8\] _1129_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__B _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4539__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__B2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6637__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4227__B1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A1 _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3838__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6214__I mod.instr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 io_in[2] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout215_I net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3530_ _3278_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3461_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__C1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ net12 _1883_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4702__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3505__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4702__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3392_ _3238_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6180_ mod.pc_1\[4\] _2869_ _2864_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _1932_ _1775_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_96_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _1208_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__B2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _0973_ _0976_ _0979_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4769__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _2421_ _2694_ _2697_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4915_ _1788_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3441__A1 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ _1812_ _1813_ _1814_ _1815_ _1805_ _1808_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_20_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ _1436_ _1746_ _1433_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3744__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ mod.registers.r15\[3\] _3095_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3728_ mod.registers.r4\[3\] _0696_ _0697_ mod.registers.r1\[3\] _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6447_ _2966_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3483__I _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3659_ mod.registers.r8\[2\] _0531_ _0532_ mod.registers.r10\[2\] _0629_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5497__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _3007_ _3000_ _3008_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5329_ mod.registers.r1\[11\] _2246_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6446__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5249__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4528__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3680__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3680__B2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4932__A1 mod.pc0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3499__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3499__B2 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4160__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__A1 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__A1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout165_I net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6802__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__S1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ _1549_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3974__A2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ mod.registers.r8\[6\] _2510_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ _1342_ _1598_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6952__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5176__B2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4562_ _0691_ _1334_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4399__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _2955_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3513_ _3217_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4493_ _1184_ _1190_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ mod.des.des_dout\[5\] _2896_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3444_ mod.registers.r11\[0\] _3292_ _0413_ mod.registers.r2\[0\] _0414_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3375_ mod.funct3\[1\] _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6163_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _1743_ _1747_ _1756_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4348__B _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout78_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _1979_ _2797_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5100__A1 mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _1178_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5651__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__I _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6996_ _0094_ net204 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5403__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5947_ mod.registers.r14\[3\] _2683_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5878_ _2554_ _2640_ _2643_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5167__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ mod.ins_ldr_3 mod.valid_out3 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_305 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_316 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_327 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_338 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_349 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6825__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3405__A1 mod.funct3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6975__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3708__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4905__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5633__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__B1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4841__C2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6850_ _0351_ net158 mod.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4615__C _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _2564_ _2591_ _2594_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _0285_ net115 mod.registers.r12\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3993_ _0485_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5732_ _2235_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5663_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _0912_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5594_ mod.registers.r6\[7\] _2454_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4545_ _1263_ _1268_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _1341_ _1054_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6215_ mod.des.des_dout\[1\] _2889_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3427_ mod.registers.r8\[0\] _3273_ _3279_ mod.registers.r10\[0\] _3280_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _2833_ _2838_ _2841_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A1 mod.registers.r1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__B2 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _1971_ _1972_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6979_ _0077_ net70 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3938__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3936__I _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5560__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4115__A2 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3874__A1 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3874__B2 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5615__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7003__CLK net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4007__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4051__A1 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout128_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4354__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _0911_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__B _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _1003_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6000_ _2711_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3865__A1 mod.registers.r15\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ _0636_ _0952_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3865__B2 mod.registers.r12\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3617__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3617__B2 mod.registers.r3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6902_ _0403_ net199 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _0334_ net187 mod.valid1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _0268_ net45 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3976_ _3241_ _0945_ _0463_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4042__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5715_ _2193_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3396__A3 mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A1 mod.registers.r10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _0199_ net55 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5646_ _2425_ _2486_ _2490_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5542__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5577_ _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6590__I0 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6670__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _1495_ _1496_ _1497_ _1432_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_104_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3491__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4459_ _1300_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6129_ mod.pc\[8\] _2048_ _1894_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3320__A3 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6307__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__C _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6022__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4033__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4497__I _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5836__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3847__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3698__I1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__I mod.instr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4960__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3830_ _0579_ _0799_ _3262_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_60_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4024__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4024__B2 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3761_ mod.registers.r8\[12\] _0729_ _0730_ mod.registers.r10\[12\] _0731_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5772__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _2161_ _2356_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3783__B1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6480_ _3077_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3692_ mod.registers.r15\[3\] _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _2236_ _2337_ _2342_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5524__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__I0 mod.des.des_dout\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _2270_ _2296_ _2297_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _1177_ _1179_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5293_ mod.registers.r1\[7\] _2206_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4244_ mod.registers.r3\[12\] _0959_ _0960_ mod.registers.r2\[12\] _0964_ mod.registers.r15\[12\]
+ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4175_ _0633_ _0712_ _1044_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout60_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4263__A1 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _0320_ net105 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4015__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__C _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4566__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _0251_ net45 mod.registers.r9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4091__B _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _0455_ _0459_ _0452_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6678_ _0182_ net58 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5629_ _2472_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6563__I0 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4006__A1 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4006__B2 mod.registers.r1\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5349__A4 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__A2 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6909__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4088__A4 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4955__I _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout195_I net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4493__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _2706_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4245__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4245__B2 mod.registers.r5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5786__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4690__I _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4862_ _3213_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _3148_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3813_ mod.registers.r7\[14\] _0743_ _0729_ mod.registers.r8\[14\] mod.registers.r12\[14\]
+ _0766_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_60_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _1741_ _1745_ _1166_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6532_ mod.registers.r15\[9\] _3107_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3744_ _0595_ _0699_ _0710_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _2147_ _3025_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3675_ mod.registers.r5\[2\] _0547_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ mod.registers.r3\[0\] _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6394_ _2123_ _2953_ _3018_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5345_ mod.des.des_dout\[34\] _2213_ _2280_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4720__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5026__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _1786_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6473__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ mod.registers.r12\[13\] _0962_ _0959_ mod.registers.r3\[13\] _0960_ mod.registers.r2\[13\]
+ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_68_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ mod.pc_2\[3\] _0778_ _1057_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__B1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3944__I mod.funct3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6161__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3514__A3 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6464__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6907__D _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4227__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4227__B2 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 mod.registers.r14\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 mod.registers.r9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3738__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 io_in[3] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ _0429_ _0410_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout208_I net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6731__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__B1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4163__C2 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3391_ _3233_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5130_ _2072_ _2073_ _2088_ _3156_ _2089_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _1909_ _1720_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6881__CLK net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ mod.registers.r13\[15\] _0980_ _0981_ mod.registers.r9\[15\] _0982_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5963_ mod.registers.r14\[9\] _2695_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4914_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3441__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4845_ mod.ldr_hzd\[3\] _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4776_ _1741_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6515_ _2396_ _3093_ _3098_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3727_ _0466_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4941__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3744__A3 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6446_ _1826_ _3047_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3658_ mod.pc_2\[2\] _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6377_ mod.pc_1\[6\] _3001_ _3004_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3589_ mod.registers.r14\[4\] _3283_ _3287_ mod.registers.r6\[4\] _0559_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5328_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3901__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _2178_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A1 mod.registers.r14\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6315__I _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6604__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5185__A2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6754__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6050__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6134__A1 mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3499__A2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__B _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout190 net191 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout158_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4620__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__B2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4630_ _1469_ _1599_ _0668_ _0924_ _0725_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4901__C mod.instr_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ _1342_ _1527_ _1530_ _1419_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6300_ _2760_ _2957_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3512_ _3183_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4492_ _1436_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6231_ mod.instr\[5\] _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3443_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4687__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _2151_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _3226_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4151__A3 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _1156_ _1160_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _2768_ _2769_ mod.pc\[4\] _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4439__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ mod.pc_2\[6\] _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5100__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6627__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3759__I _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6995_ _0093_ net209 mod.des.des_dout\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__I _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ _2396_ _2681_ _2686_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ mod.registers.r12\[9\] _2641_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _1191_ _0907_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5167__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__A1 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ _1538_ _1301_ _1537_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_5_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3494__I _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ _3029_ _3041_ _3038_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3350__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A2 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_306 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_317 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_328 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_339 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3405__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5884__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6355__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6107__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A1 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5330__A2 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4841__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__B2 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5800_ mod.registers.r10\[13\] _2592_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6780_ _0284_ net77 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3992_ _0888_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _2546_ _2541_ _2547_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6830__D _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6346__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _1071_ _1452_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _2411_ _2453_ _2457_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4544_ _1269_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3580__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4109__B1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1072_ _1063_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ mod.instr\[1\] _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3426_ _3278_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _2833_ _2838_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _3209_ _3187_ _3206_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5034__I mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _2781_ _1913_ _1797_ _2770_ _2775_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5969__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5027_ mod.pc_2\[4\] _1972_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6978_ _0076_ net69 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _2430_ _2673_ _2675_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__C _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5209__I _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A1 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3874__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5076__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6942__CLK net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3399__I _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3929__A3 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4051__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5000__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _1227_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5282__C _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4191_ _1152_ _1156_ _1160_ _1143_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3865__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5067__A1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__B _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3617__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6901_ _0402_ net198 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6832_ _0333_ net186 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6763_ _0267_ net45 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3975_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5714_ _2534_ _2530_ _2535_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _0198_ net57 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ mod.registers.r7\[10\] _2487_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _2444_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6590__I1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _1492_ _1444_ _1456_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4458_ _1296_ _3242_ _1399_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3409_ _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4389_ _1356_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6128_ mod.pc\[9\] _2065_ _1894_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4817__B _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ _2764_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4552__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4033__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__A1 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__I0 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3847__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3480__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4024__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6838__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _0500_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__A1 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3783__B2 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ _0417_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5430_ mod.registers.r3\[7\] _2338_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5524__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__B _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6988__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ mod.registers.r1\[15\] _2277_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _1279_ _1280_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5288__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _1209_ _1210_ _1211_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4174_ _0595_ _1131_ _1142_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout53_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5460__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _0319_ net101 mod.registers.r14\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6746_ _0250_ net49 mod.registers.r9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3958_ _0925_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4566__A3 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3369__A4 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3774__A1 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3889_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6677_ _0181_ net57 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5982__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _2400_ _2473_ _2479_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6563__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__I0 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5559_ mod.registers.r5\[12\] _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4547__B _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3462__B1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4006__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__B1 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6554__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5690__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout188_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6660__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4930_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5288__B _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3587__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4861_ _1781_ _1191_ _0907_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6600_ net7 mod.des.des_dout\[35\] _3136_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3812_ mod.registers.r3\[14\] _0752_ _0736_ mod.registers.r2\[14\] _0782_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _1436_ _1760_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5745__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6531_ _2416_ _3106_ _3108_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3743_ _0615_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6462_ _1817_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3674_ mod.registers.r7\[2\] _0548_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5413_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6393_ mod.pc_1\[12\] _2720_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5344_ _2166_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5275_ _2171_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _1192_ _1193_ _1194_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5130__B1 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4157_ _1125_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _0657_ _0658_ _0659_ _0664_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3698__S _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3444__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__A1 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3995__B2 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6729_ _0233_ net46 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5217__I _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3514__A4 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5672__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3683__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4227__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A1 mod.registers.r3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3435__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3738__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3738__B2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__B _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 io_in[4] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4163__A1 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout103_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__B2 mod.registers.r4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3390_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4966__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3910__A1 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3870__I _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _2021_ _2022_ _2023_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ _0603_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _2416_ _2694_ _2696_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5966__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3977__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ _1801_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5893_ _2161_ _2624_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__B1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ mod.ldr_hzd\[2\] _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4775_ _1188_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6391__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6514_ mod.registers.r15\[2\] _3095_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3726_ _0465_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _3052_ _3053_ _3046_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3657_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6143__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3588_ mod.registers.r7\[4\] _0442_ _3273_ mod.registers.r8\[4\] _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6376_ _2008_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3901__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3901__B2 mod.registers.r7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5327_ mod.des.des_dout\[32\] _2248_ _2264_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_130_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5654__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4209_ _3239_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5189_ _2140_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5406__A1 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4209__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4145__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__C _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4448__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5645__A1 mod.registers.r7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout180 net181 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout191 net193 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A3 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4454__C _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__A1 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4560_ _0811_ _1528_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3511_ _0480_ _3256_ mod.registers.r14\[1\] _0477_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4491_ _1459_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _2903_ _2901_ _2904_ _2905_ _2898_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3442_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3373_ mod.funct3\[2\] _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6161_ _2131_ _2824_ _2853_ _2854_ _2855_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _1962_ _2766_ _2796_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4439__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1932_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__B _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5320__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _0092_ net209 mod.des.des_dout\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5945_ mod.registers.r14\[2\] _2683_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5876_ _2550_ _2640_ _2642_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _1389_ _1788_ _1791_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__3775__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4375__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4758_ _1724_ _1384_ _1725_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3709_ _0675_ _0676_ _0677_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5990__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ _0942_ _0914_ _0915_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _1858_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5875__A1 mod.registers.r12\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__B mod.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6359_ _2872_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3886__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_307 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_318 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_329 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__I _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6052__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6061__I _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4366__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6871__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__A2 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5866__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3341__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout170_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ mod.registers.r3\[15\] _0959_ _0960_ mod.registers.r2\[15\] _0961_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5730_ mod.registers.r9\[6\] _2542_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5661_ _2357_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4612_ _1580_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5592_ mod.registers.r6\[6\] _2454_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _1512_ _1439_ _1438_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4109__A1 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__B2 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _1437_ _1256_ _1441_ _1443_ _1257_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__A1 mod.registers.r12\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6213_ _2887_ _2719_ _2890_ _2892_ _2855_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3425_ _3267_ _3269_ _3275_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout83_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6144_ _2101_ _2840_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3356_ _3158_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ mod.pc\[1\] _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _1163_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6744__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6977_ _0075_ net123 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6894__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ mod.registers.r13\[12\] _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3719__B _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ mod.registers.r12\[2\] _2629_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4348__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5848__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3859__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5076__A2 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__B1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5895__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__B _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4339__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5000__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6617__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4190_ _1157_ _1158_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5067__A2 _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _0401_ net166 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4814__B3 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _0002_ _0006_ net206 mod.des.des_counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__4027__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _0266_ net81 mod.registers.r10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _0942_ _0943_ _0915_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4042__A3 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5713_ mod.registers.r9\[1\] _2532_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3539__B _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ _0197_ net57 mod.registers.r6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5644_ _2422_ _2486_ _2489_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5575_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4526_ _1259_ _1271_ _1151_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4750__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4457_ _1418_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5045__I _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3408_ _3253_ _3180_ _3222_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4388_ _1357_ _0840_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _2817_ _2820_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ mod.registers.r6\[0\] _3186_ _3189_ mod.registers.r5\[0\] mod.registers.r2\[0\]
+ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_85_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _1953_ _1973_ _1954_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__B _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__A2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3792__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4344__I1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5049__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4009__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3480__A1 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3480__B2 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5221__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout133_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ mod.registers.r12\[3\] _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__I mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4311_ _0874_ _1121_ _1123_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ mod.des.des_dout\[28\] _2188_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5288__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4242_ mod.registers.r12\[12\] _0962_ _0975_ mod.registers.r1\[12\] _1212_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _1021_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4799__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5460__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout46_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6814_ _0318_ net105 mod.registers.r14\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _0249_ net48 mod.registers.r9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3957_ _0926_ _0774_ _0453_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3774__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _0180_ net103 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3888_ _0843_ _3239_ _0852_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4879__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5627_ mod.registers.r7\[3\] _2475_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6932__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4184__C1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4574__I1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _2390_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _1329_ _1472_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5489_ _2361_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5279__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4119__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5451__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3462__A1 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3462__B2 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5203__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4714__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6805__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__I1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4860_ _1803_ _1811_ _1829_ _3244_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3811_ mod.registers.r15\[14\] _0765_ _0751_ mod.registers.r9\[14\] _0781_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _1273_ _1278_ _1759_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ mod.registers.r15\[8\] _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3742_ mod.funct7\[0\] _0711_ _0617_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4699__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _3032_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3673_ _0629_ _0630_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4705__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ _2328_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6392_ _2752_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _2042_ _2241_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _2201_ _2218_ _2219_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4225_ mod.registers.r1\[13\] _0975_ _0981_ mod.registers.r9\[13\] _1195_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5130__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4156_ _0873_ _1124_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4087_ _0652_ _0653_ _0654_ _0655_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3778__I mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__B _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3444__B2 mod.registers.r2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _1952_ _1955_ _1794_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6728_ _0232_ net54 mod.registers.r8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _0163_ net146 mod.registers.r4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__B _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3683__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3683__B2 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6978__CLK net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3435__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3435__B2 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3738__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4935__B2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput15 io_in[5] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _0608_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3674__A1 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ mod.registers.r14\[8\] _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4912_ _1830_ _1876_ _1881_ _1817_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3977__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5892_ _2568_ _2646_ _2651_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5179__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ mod.ldr_hzd\[1\] _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4774_ _1102_ _1105_ _1279_ _1492_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _2393_ _3093_ _3097_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3725_ mod.registers.r3\[3\] _0694_ _0596_ mod.registers.r7\[3\] _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _2967_ _3041_ _3037_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3656_ _0625_ _0622_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4154__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5351__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _0580_ _3000_ _3006_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3587_ _0459_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5326_ _2166_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3901__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ mod.des.des_dout\[25\] _2167_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5053__I mod.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ _0424_ _0953_ _0956_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5188_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _1107_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5406__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3301__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4090__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A1 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5228__I _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5342__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4145__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5893__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4288__B _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__I _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5645__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7006__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout170 net171 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3656__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout181 net201 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout192 net193 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3671__A4 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__B1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3959__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5581__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout213_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3510_ _3209_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4490_ _1224_ _1276_ _1286_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5333__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3441_ _3275_ _3277_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _2788_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3372_ _3154_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A1 mod.registers.r11\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__B2 mod.registers.r2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5111_ _0000_ mod.des.des_counter\[1\] _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _0003_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5042_ _1685_ _1696_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__C _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6993_ _0091_ net212 mod.des.des_dout\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _2393_ _2681_ _2685_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ mod.registers.r12\[8\] _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6432__I _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4826_ _1794_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _1699_ _1723_ _1726_ _1247_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6673__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ mod.registers.r9\[1\] _0511_ _0500_ mod.registers.r10\[1\] _0678_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4688_ _1383_ _1650_ _1653_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5324__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _1814_ _3033_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3639_ mod.registers.r12\[2\] _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6358_ _2952_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3886__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5309_ _1972_ _2241_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3350__A3 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ mod.des.des_dout\[20\] _2900_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_308 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_319 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5511__I _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__I0 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__A2 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A1 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6342__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4366__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3326__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__A2 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A2 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _0701_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__B _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _2146_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4611_ _1267_ _1264_ _1266_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5554__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5591_ _2408_ _2453_ _2456_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _1448_ _1453_ _1454_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4109__A2 _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _1097_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6212_ _2891_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5857__A2 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3424_ _3276_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_98_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ mod.pc\[11\] _1914_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3355_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout76_I net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6074_ _2765_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5025_ _1082_ _1087_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6034__A2 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6976_ _0074_ net122 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5927_ _2655_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5793__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _2534_ _2627_ _2631_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4809_ _1390_ _1394_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5545__A1 mod.registers.r5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5789_ _2550_ _2585_ _2587_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3859__A1 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4520__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6337__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4036__A1 mod.registers.r2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__B2 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 mod.registers.r10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4511__A2 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _0001_ _0005_ net206 mod.des.des_counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XANTENNA__4027__A1 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4027__B2 mod.registers.r5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6761_ _0265_ net81 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5775__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3973_ _0935_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _2185_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4042__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6692_ _0196_ net103 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5643_ mod.registers.r7\[9\] _2487_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5527__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4525_ _0912_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _1235_ _1371_ _1424_ _1331_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6711__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3407_ _3254_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4502__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _0460_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ mod.pc\[9\] _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4266__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ mod.pc_2\[3\] _1951_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5996__I _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4018__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4833__C _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _0057_ net216 mod.des.des_dout\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5518__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__I _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4140__I _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3701__B1 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6067__I _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4257__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4009__A1 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__B2 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3480__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4980__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout126_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4310_ _0859_ _1144_ _1146_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5290_ _2231_ _2232_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4241_ mod.registers.r14\[12\] _0977_ _0978_ mod.registers.r7\[12\] _1211_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4172_ _1132_ _1133_ _1140_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_68_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4799__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5748__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _0317_ net101 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout39_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6744_ _0248_ net64 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3956_ _3246_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6675_ _0179_ net104 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3887_ _0853_ _0854_ _0855_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5626_ _2397_ _2473_ _2478_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6173__A1 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4184__B1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _2388_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4184__C2 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__A1 mod.registers.r13\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4508_ _1473_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _2359_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4439_ _0757_ _0774_ _1291_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _2808_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4239__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__B2 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3462__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4411__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4962__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5911__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3922__B1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A1 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3453__A2 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3810_ mod.registers.r5\[14\] _0741_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _1278_ _1759_ _1273_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _3215_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _2716_ _3063_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3672_ _0498_ _0635_ _0639_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5411_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4705__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6391_ _2095_ _2953_ _3016_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5902__A1 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5342_ _0758_ _2181_ _2214_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3913__B1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4929__B _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3833__B _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5273_ mod.registers.r1\[5\] _2206_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4469__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ mod.registers.r14\[13\] _0977_ _0889_ mod.registers.r13\[13\] _0978_ mod.registers.r7\[13\]
+ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5130__A2 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4155_ _0873_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3444__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _1953_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6727_ _0231_ net54 mod.registers.r8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3939_ mod.funct7\[1\] _0905_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _0162_ net146 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _2431_ _2465_ _2467_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6589_ _3135_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4172__A3 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3683__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4632__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3435__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 io_in[6] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6137__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3371__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout193_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3674__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6255__I mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5960_ _2682_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4911_ _1877_ _1878_ _1879_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5891_ mod.registers.r12\[15\] _2647_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ mod.ldr_hzd\[0\] _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ _1740_ _1742_ _1699_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6604__RN _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3724_ _0471_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6512_ mod.registers.r15\[1\] _3095_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _1822_ _3047_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3655_ _0495_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6374_ mod.pc_1\[5\] _3001_ _3004_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3586_ _0455_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5325_ _2009_ _2241_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5334__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _2181_ _1968_ _2173_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6300__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _1152_ _1171_ _1176_ _1143_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_102_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ net11 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3665__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ mod.registers.r3\[9\] _0694_ _0882_ mod.registers.r5\[9\] _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3789__I _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__I _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input19_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4069_ mod.registers.r1\[6\] _0466_ _3204_ mod.registers.r8\[6\] _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4614__A1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3417__A2 mod.instr_2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4090__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4413__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A3 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6945__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout160 net161 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout171 net173 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4853__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout182 net188 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout193 net194 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3699__I mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__I mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3408__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__B2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3959__A3 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3813__C1 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__A3 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3440_ _3284_ _3268_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_fanout206_I net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6530__A1 mod.registers.r15\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3371_ _3180_ _3222_ _3223_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _1908_ _2055_ _2069_ _0001_ _2070_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__3895__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _2792_ _2794_ _2773_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5041_ _1916_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3402__I mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ _0090_ net210 mod.des.des_dout\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5943_ mod.registers.r14\[1\] _2683_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5874_ _2628_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ mod.pc_2\[0\] _1078_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5021__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5572__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _1724_ _1725_ _1302_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3707_ mod.registers.r5\[1\] _0517_ _0518_ mod.registers.r7\[1\] _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _1243_ _1655_ _1656_ _1433_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3638_ _3210_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6426_ _3035_ _3039_ _3023_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6521__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6968__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3335__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6357_ _2992_ _2994_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3569_ _0533_ _0536_ _0537_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3886__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5308_ _2191_ _2055_ _2209_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ mod.instr\[20\] _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_309 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _2165_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__I _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__I1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 mod.registers.r1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3810__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5239__I _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5563__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6512__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__B2 mod.registers.r1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3629__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout156_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _1449_ _1451_ _1452_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5590_ mod.registers.r6\[5\] _2454_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4541_ _1494_ _1498_ _1499_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4762__B1 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3892__I mod.pc_2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4472_ _1048_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6211_ net13 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3423_ mod.instr_2\[10\] _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _2832_ _2839_ _2831_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3354_ _3183_ _3184_ _3206_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _2774_ _2777_ _2779_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1987_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout69_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A1 mod.registers.r4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__B _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6975_ _0073_ net122 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ _2653_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6640__CLK net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5793__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5857_ mod.registers.r12\[1\] _2629_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4808_ _1376_ _1698_ _1758_ _1775_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5545__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ mod.registers.r10\[8\] _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6790__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _1635_ _1636_ _1343_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _1850_ _2883_ _3027_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5522__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A1 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6554__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__B _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__A1 mod.pc_2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4036__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6353__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5536__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6528__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5472__A1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4275__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6663__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4027__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5224__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__I mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6760_ _0264_ net65 mod.registers.r10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _3248_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _2527_ _2530_ _2533_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ _0195_ net103 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5642_ _2417_ _2486_ _2488_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ _2299_ _2356_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5607__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4524_ _1491_ _1493_ _1242_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4455_ _1004_ _0934_ _1246_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ _3255_ _3256_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4386_ _0813_ _0814_ _0826_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3710__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3710__B2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6125_ _2818_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3337_ _3182_ _3159_ _3163_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6056_ _2725_ _1899_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_85_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4266__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ mod.pc_2\[3\] _1951_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A2 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _0056_ net215 mod.des.des_dout\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5909_ _2402_ _2661_ _2663_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6889_ _0390_ net170 mod.instr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4726__B1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4421__I _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6348__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3701__A1 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3701__B2 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6686__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5206__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6083__I _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4331__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3940__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ mod.registers.r11\[12\] _0974_ _0980_ mod.registers.r13\[12\] _1210_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5693__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4171_ mod.registers.r2\[8\] _0893_ _0468_ mod.registers.r5\[8\] mod.registers.r11\[8\]
+ _0605_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A1 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6812_ _0316_ net44 mod.registers.r13\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5748__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6743_ _0247_ net66 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3955_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6674_ _0178_ net104 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3886_ mod.registers.r5\[8\] _0440_ _0413_ mod.registers.r2\[8\] _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5625_ mod.registers.r7\[2\] _2475_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5337__I _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4184__A1 mod.registers.r5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4184__B2 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5556_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5920__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4507_ _0811_ _1474_ _1475_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5487_ _2268_ _2373_ _2378_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _1404_ _1407_ _1351_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4369_ _1336_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _2016_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4239__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__A1 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6039_ _2139_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5021__B _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5739__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6400__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4411__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3922__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3922__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3990__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5427__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__B _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4402__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _0702_ _0704_ _0707_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5157__I mod.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ _0637_ _0445_ mod.registers.r2\[2\] _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5410_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ mod.pc_1\[11\] _2720_ _3012_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4996__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3913__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5341_ _2182_ _2122_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3913__B2 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5272_ _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4469__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__A1 mod.registers.r8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ mod.registers.r6\[13\] _0966_ _0967_ mod.registers.r5\[13\] _1193_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3677__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4154_ _1121_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4437__S _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4085_ _0759_ _0620_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5620__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4680__B _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _1051_ _1935_ _1917_ _1937_ _1938_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6394__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__I _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _0230_ net59 mod.registers.r8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3938_ _0902_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3601__B1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ _0161_ net136 mod.registers.r4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3869_ mod.pc_2\[10\] _0778_ _0833_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5608_ mod.registers.r6\[12\] _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6588_ _3141_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5539_ _2388_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5657__A1 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5530__I _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3985__I mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6874__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 io_in[7] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6137__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3371__A2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5648__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout186_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6073__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4910_ _1815_ _1814_ _1813_ _1812_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5890_ _2566_ _2646_ _2650_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _1804_ _1806_ _0661_ _1807_ _1809_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_33_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__I mod.instr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _1741_ _1281_ _1650_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6511_ _2385_ _3093_ _3096_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3723_ _0627_ _0668_ _0686_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _3050_ _3051_ _3046_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3654_ _0497_ _0555_ _0594_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5887__A1 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6373_ _3003_ _3000_ _3005_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3585_ _0526_ _0527_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3898__B1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ _2191_ _2090_ _2214_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout99_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5255_ _1971_ _2182_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4311__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _1172_ _1173_ _1174_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_68_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6747__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5186_ _2138_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3665__A3 mod.registers.r11\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ mod.registers.r10\[9\] _1106_ _0703_ mod.registers.r9\[9\] _1107_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6064__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ mod.registers.r3\[6\] _0471_ _0465_ mod.registers.r4\[6\] _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5811__A1 mod.registers.r11\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6897__CLK net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__B1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _0213_ net61 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__A1 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5525__I _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4145__A4 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3353__A2 mod.instr_2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4302__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_94_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout161 net162 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout172 net173 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout183 net188 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout194 net200 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6055__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__A1 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3408__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__B1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__C2 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6602__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4369__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A3 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5030__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5869__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout101_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3370_ _3153_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5097__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _1787_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__B _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6266__I mod.instr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6046__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6991_ _0089_ net212 mod.des.des_dout\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _2385_ _2681_ _2684_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5873_ _2626_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4514__I _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _1792_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5021__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _1204_ _1459_ _1292_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4780__A1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3706_ mod.registers.r14\[1\] _0502_ _3291_ mod.registers.r11\[1\] _0676_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ _1506_ _1493_ _1651_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6425_ _3029_ _3036_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3637_ _3207_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6356_ _0955_ _2989_ _2962_ mod.instr\[20\] _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3568_ mod.registers.r4\[7\] _0508_ _3237_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ mod.pc_2\[9\] _2221_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6287_ _2946_ _2889_ _2947_ _2941_ _2742_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3499_ mod.registers.r2\[1\] _3191_ _0468_ mod.registers.r5\[1\] _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _2164_ _2186_ _2187_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4296__B1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _2124_ _2111_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4424__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4523__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3326__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3877__A3 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3503__I _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__B1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4540_ _1504_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _1438_ _1439_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6210_ mod.des.des_dout\[0\] _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3422_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2834_ _2836_ _2838_ _2817_ _2773_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_97_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3353_ _3161_ mod.instr_2\[16\] _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ mod.pc\[1\] _2774_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5114__B _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _3243_ _1554_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3413__I _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6019__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _0072_ net125 mod.registers.r15\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ _2427_ _2667_ _2672_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5856_ _2527_ _2627_ _2630_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4807_ _1392_ _1395_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6935__CLK net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4202__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5787_ _2573_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4738_ _1429_ _0901_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4669_ _0717_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ mod.rd_3\[0\] _2884_ _3017_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _2978_ _2983_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4419__I _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5481__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__B _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3993__I _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__C _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6808__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__B _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5224__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6421__A1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__CLK net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3971_ _0929_ _0934_ _0685_ _0938_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ mod.registers.r9\[0\] _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4983__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6690_ _0194_ net103 mod.registers.r6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ mod.registers.r7\[8\] _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5572_ _2442_ _2432_ _2443_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1102_ _1105_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5109__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ _1420_ _1421_ _1423_ _1340_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3405_ mod.funct3\[2\] _3232_ _3257_ _3234_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _1353_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout81_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _2050_ _2780_ _2823_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3710__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3336_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _2734_ _2134_ _2763_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5006_ _1122_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _0055_ net215 mod.des.des_dout\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5908_ mod.registers.r13\[4\] _2662_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6888_ _0389_ net170 mod.instr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _2598_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__B2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5151__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4593__B _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__B1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__I _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__A1 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5443__I _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6630__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _1134_ _1137_ _1138_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6780__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _0315_ net48 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _0246_ net70 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3954_ _0923_ _0808_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ _0177_ net99 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3885_ mod.registers.r14\[8\] _3283_ _0428_ mod.registers.r9\[8\] _0855_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4708__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5624_ _2394_ _2473_ _2477_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5381__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ _2275_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4184__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4506_ _1316_ _0927_ _1350_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ mod.registers.r4\[11\] _2374_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6449__I _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _1405_ _0462_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5353__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4368_ _1337_ _0724_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _2802_ _1885_ mod.pc\[6\] _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3319_ _3158_ _3159_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0899_ _1251_ _1075_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6038_ _2730_ _2053_ _2751_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6184__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5021__C _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A4 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__C _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5372__A1 mod.registers.r2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3922__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5124__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__I _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3686__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ _0631_ _0562_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5363__A1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ _2270_ _2276_ _2278_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__I _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ mod.des.des_dout\[26\] _2188_ _2212_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_4222_ mod.registers.r15\[13\] _0964_ _0968_ mod.registers.r8\[13\] _1192_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3677__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3677__B2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4153_ _0577_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _1051_ _0499_ _1052_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__3429__A1 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_290 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4641__A3 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout44_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _1051_ _1935_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6725_ _0229_ net61 mod.registers.r8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3937_ _0904_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3601__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3601__B2 mod.registers.r11\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _0160_ net131 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3868_ _0834_ _0835_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_109_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _2447_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5354__A1 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ net19 mod.des.des_dout\[29\] _3137_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3799_ mod.registers.r9\[13\] _0428_ _0752_ mod.registers.r3\[13\] _0769_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5469_ _2361_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3668__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5409__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4396__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5258__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 io_in[8] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5345__A1 mod.des.des_dout\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__A1 mod.registers.r8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3659__B2 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4337__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4084__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout179_I net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4084__B2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6699__CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ mod.ldr_hzd\[10\] _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4771_ _1272_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5584__A1 mod.registers.r6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ mod.registers.r15\[0\] _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3722_ _0691_ _0622_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3595__B1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6441_ _2967_ _3036_ _3037_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5336__A1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3653_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3347__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ mod.pc_1\[4\] _3001_ _3004_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3584_ _0529_ _0551_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_127_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3898__A1 mod.registers.r15\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5323_ mod.pc_2\[11\] _2169_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5254_ _2163_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ mod.registers.r12\[11\] _1110_ _0882_ mod.registers.r5\[11\] _0696_ mod.registers.r4\[11\]
+ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4311__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ _1781_ net22 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _3195_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A2 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4067_ _1034_ _1035_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4075__A1 mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3822__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__B2 mod.registers.r7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4969_ _0954_ _0492_ _1936_ _0669_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_51_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _0212_ net106 mod.registers.r7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__A1 mod.des.des_dout\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6639_ _0143_ net129 mod.registers.r3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4302__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout151 net152 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout162 net202 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout173 net180 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout184 net187 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout195 net197 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__A1 mod.registers.r5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__B2 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__A1 mod.registers.r7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3996__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3813__B2 mod.registers.r8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6602__I1 mod.des.des_dout\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__CLK net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6483__S _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4057__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _0088_ net210 mod.des.des_dout\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5941_ mod.registers.r14\[0\] _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ _2548_ _2634_ _2639_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4823_ _0903_ _0906_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _1287_ _1293_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5309__A1 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3705_ mod.registers.r15\[1\] _0514_ _0512_ mod.registers.r3\[1\] _0675_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _1651_ _1506_ _1493_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4780__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6424_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3636_ mod.registers.r11\[2\] _0605_ _0473_ mod.registers.r8\[2\] _0606_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _2992_ _2993_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3567_ mod.registers.r11\[7\] _0505_ _0506_ mod.registers.r2\[7\] _0537_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3335__A3 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5306_ _2165_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6286_ mod.des.des_dout\[19\] _2900_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3498_ _3188_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5237_ mod.registers.r1\[1\] _2179_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4296__B2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _2123_ _1089_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4119_ mod.funct7\[2\] _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ mod.pc_2\[9\] _1233_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6596__I0 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4220__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4523__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6568__S _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A2 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4039__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4039__B2 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__B1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6587__I0 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4211__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4762__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout211_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _1253_ _1099_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3421_ mod.instr_2\[11\] _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5711__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3352_ mod.registers.r11\[0\] _3202_ _3204_ mod.registers.r8\[0\] _3205_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6277__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _2753_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4278__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _3154_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _0071_ net114 mod.registers.r15\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5924_ mod.registers.r13\[11\] _2668_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5855_ mod.registers.r12\[0\] _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _1394_ _1698_ _1758_ _1775_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4202__A1 mod.registers.r3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4202__B2 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _2571_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4753__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _1701_ _1702_ _1384_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4668_ _0811_ _1635_ _1636_ _1637_ _1468_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4505__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _3025_ _3026_ _3023_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3619_ mod.registers.r13\[5\] _0446_ _0448_ mod.registers.r1\[5\] _0589_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _0809_ _1532_ _1534_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ _0846_ _2982_ _2979_ mod.instr\[13\] _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6258__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _2741_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A3 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3492__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5769__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A2 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4744__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5941__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__I _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout161_I net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4432__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4983__A2 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5640_ _2474_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5571_ mod.registers.r5\[15\] _2433_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5932__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4522_ _1490_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3943__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4453_ _1242_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4948__C _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3404_ mod.instr_2\[2\] mod.instr_2\[0\] _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4384_ _0683_ _0684_ _0859_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6123_ _2765_ _2821_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3335_ _3166_ _3167_ _3175_ _3187_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ mod.pc0\[13\] _2723_ _2754_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5999__A1 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ mod.pc_2\[4\] _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6902__CLK net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _0054_ net196 mod.ldr_hzd\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4423__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5907_ _2655_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4974__A2 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6887_ _0388_ net171 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__C1 mod.registers.r2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6176__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ _2558_ _2612_ _2617_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__B1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _2527_ _2572_ _2575_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__B _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__A3 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__B2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__A2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6581__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4965__A2 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4717__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__A1 mod.registers.r13\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__CLK net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6810_ _0314_ net66 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6741_ _0245_ net69 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3953_ _0625_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3884_ mod.registers.r13\[8\] _0447_ _3279_ mod.registers.r10\[8\] _0854_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _0176_ net58 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5623_ mod.registers.r7\[1\] _2475_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5905__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3419__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5554_ _2428_ _2418_ _2429_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _1401_ _1310_ _0575_ _0812_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5485_ _2261_ _2373_ _2377_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4436_ _0801_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ _1250_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _2783_ _2791_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3318_ mod.registers.r3\[0\] _3165_ _3170_ mod.registers.r7\[0\] _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _1264_ _1266_ _1267_ _1260_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6037_ _2729_ mod.pc0\[8\] _2731_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4644__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4644__B2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6939_ _0037_ net195 mod.rd_3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6149__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3329__I mod.instr_2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__B _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__CLK net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6576__S _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3686__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4635__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6388__A1 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5270_ _2213_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ _0720_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3677__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4874__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4152_ _0637_ _0897_ _1044_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__B1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _0644_ _0645_ _0646_ _0648_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3429__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_280 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_291 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5051__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _0651_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5629__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _0228_ net106 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3601__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _0159_ net133 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3867_ mod.registers.r13\[10\] _0745_ _0746_ mod.registers.r1\[10\] _0837_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5606_ _2445_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5354__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6586_ _3140_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3798_ mod.registers.r13\[13\] _0447_ _0449_ mod.registers.r1\[13\] _0768_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3365__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5537_ _2244_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _2359_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ _2303_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3668__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4865__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6620__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5593__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 io_in[9] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6542__A1 mod.registers.r15\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3659__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3522__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__C1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4084__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__B _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _1738_ _1739_ _1167_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3721_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ _1824_ _3047_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3652_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3347__B2 mod.registers.r9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3583_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6371_ _2872_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3898__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ _2238_ _2261_ _2262_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _2164_ _2199_ _2200_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ mod.registers.r8\[11\] _0706_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5184_ _2137_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4311__A3 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _1031_ _0525_ _1103_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_29_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ mod.registers.r5\[6\] _3189_ _3199_ mod.registers.r9\[6\] _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _3229_ _0954_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6793__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6707_ _0211_ net120 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _3211_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4899_ _1861_ _1867_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6638_ _0142_ net129 mod.registers.r3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6524__A1 mod.registers.r15\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3607__I _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _3130_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout130 net132 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout141 net149 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout152 net203 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout163 net167 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout174 net175 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3342__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout185 net187 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout196 net197 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4066__A2 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3813__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5015__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__I _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout191_I net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6666__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5871_ mod.registers.r12\[7\] _2635_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4822_ _1191_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3568__A1 mod.registers.r4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__B1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4753_ _1722_ _1204_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5907__I _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _0670_ _0671_ _0672_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4684_ _1650_ _1653_ _1429_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6423_ mod.instr_2\[6\] _3025_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3635_ _3201_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6354_ mod.funct7\[1\] _2989_ _2962_ mod.instr\[19\] _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3566_ mod.registers.r14\[7\] _0534_ _0535_ mod.registers.r6\[7\] _0536_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3871__B _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _2238_ _2245_ _2247_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ mod.instr\[19\] _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3497_ mod.registers.r4\[1\] _0465_ _0466_ mod.registers.r1\[1\] _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5236_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _2123_ _1089_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4118_ _1082_ _1087_ _0457_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5098_ _2057_ _2045_ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input17_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4049_ mod.registers.r14\[7\] _0607_ _0596_ mod.registers.r7\[7\] _1019_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4205__C1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6596__I1 mod.des.des_dout\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__S0 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6141__C _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__B1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__I _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6689__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5484__A1 mod.registers.r4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4039__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3798__A1 mod.registers.r13\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3798__B2 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6587__I1 mod.des.des_dout\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4211__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3420_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3722__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__I _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3351_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _2771_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ _1908_ _1968_ _1984_ _1986_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _0070_ net114 mod.registers.r15\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5923_ _2424_ _2667_ _2671_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ _2628_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4805_ _1762_ _1765_ _1766_ _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5785_ _2548_ _2579_ _2584_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4202__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _1699_ _1701_ _1702_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4667_ _1350_ _1334_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__CLK net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ mod.ins_ldr_3 _2995_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3618_ mod.registers.r5\[5\] _0439_ _0441_ mod.registers.r7\[5\] _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5702__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__B _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _1524_ _1526_ _0623_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6337_ _2860_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3549_ mod.registers.r5\[6\] _0517_ _0518_ mod.registers.r7\[6\] _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6268_ mod.des.des_dout\[14\] _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4269__A2 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5466__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A4 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5219_ _2169_ _1387_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ mod.pc_1\[11\] _2877_ _2880_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4992__A3 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5547__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__B1 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3468__B1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3530__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4432__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout154_I net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6854__CLK net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2441_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5932__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4521_ _1102_ _1105_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3943__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3943__B2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4452_ _0923_ _1305_ _0950_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__I mod.instr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3403_ _3187_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _0926_ _0774_ _0874_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5192__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _2753_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3334_ _3176_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5448__A1 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _2760_ _2762_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _1794_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout67_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4671__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__I _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _0053_ net196 mod.ldr_hzd\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5906_ _2653_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6886_ _0387_ net171 mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__B1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3631__C2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ mod.registers.r11\[11\] _2613_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5367__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6176__A2 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__A1 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4187__B2 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ mod.registers.r10\[0\] _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1307_ _1598_ _1688_ _1328_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_163_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _2436_ _2521_ _2524_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5687__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5439__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5830__I _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4874__C _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4111__A1 mod.registers.r5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4111__B2 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6147__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6877__CLK net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4178__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4717__A3 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5678__A1 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4130__B _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3689__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4350__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__C _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__A2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5602__A1 mod.registers.r6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _0244_ net125 mod.registers.r9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3613__B1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6671_ _0175_ net98 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5187__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3883_ mod.registers.r1\[8\] _0449_ _0431_ mod.registers.r3\[8\] _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6158__A2 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__A1 mod.registers.r3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _2386_ _2473_ _2476_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ mod.registers.r5\[11\] _2419_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _0461_ _1054_ _0682_ _0923_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5484_ mod.registers.r4\[10\] _2374_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _0461_ _1054_ _0682_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4341__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4366_ _0878_ _1241_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _1979_ _2797_ _1998_ _2803_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3317_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5650__I _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _1055_ _1061_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2743_ _2750_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5841__A1 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _0036_ net195 mod.rd_3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _0370_ net192 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3907__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6430__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4635__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6592__S _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5735__I _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _1180_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4795__B _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3677__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4874__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _3253_ _1109_ _1120_ _1021_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_110_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6076__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4082_ _0629_ _0630_ _0642_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3429__A3 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A1 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_270 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_281 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_292 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _1145_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5051__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6723_ _0227_ net122 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3935_ _3231_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6654_ _0158_ net132 mod.registers.r4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3866_ mod.registers.r5\[10\] _0741_ _0743_ mod.registers.r7\[10\] _0836_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5605_ _2428_ _2459_ _2464_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6585_ net18 mod.des.des_dout\[28\] _3137_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3797_ mod.registers.r15\[13\] _0765_ _0766_ mod.registers.r12\[13\] _0767_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4562__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _2414_ _2404_ _2415_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5467_ _2199_ _2360_ _2366_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4418_ mod.valid2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5398_ _2301_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4865__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6476__I _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4349_ _1074_ _0527_ _0573_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4617__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6019_ _2734_ mod.pc0\[3\] _2737_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3825__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__I _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6542__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3803__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4069__B1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__B1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__C2 mod.registers.r6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3678__C _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6230__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__B1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3720_ _0688_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4792__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3595__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3651_ _0578_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6533__A2 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3347__A2 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1971_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3582_ _3261_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5321_ mod.registers.r1\[10\] _2246_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6497__S _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ mod.registers.r1\[3\] _2179_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ mod.registers.r15\[11\] _0884_ _1106_ mod.registers.r10\[11\] _1173_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3713__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5183_ _1792_ _0907_ _1887_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _1030_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4065_ mod.registers.r15\[6\] _0963_ _3186_ mod.registers.r6\[6\] _1035_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4967_ _1025_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3918_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6706_ _0210_ net120 mod.registers.r7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4898_ mod.ldr_hzd\[14\] _1857_ _1853_ mod.ldr_hzd\[13\] mod.ldr_hzd\[12\] _1856_
+ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6637_ _0141_ net93 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3849_ _0815_ _0816_ _0817_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ mod.des.des_dout\[21\] net6 _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _2204_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ mod.des.des_dout\[10\] net8 _3085_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout120 net121 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3623__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout142 net144 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout153 net155 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout164 net167 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout175 net179 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout186 net187 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout197 net198 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6460__A1 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__B1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4390__S _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4774__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4526__A1 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3533__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout184_I net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4057__A3 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _2546_ _2634_ _2638_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _1790_ _1387_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3568__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _1222_ _1463_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4765__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__B2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ mod.registers.r4\[1\] _0419_ _3264_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _1651_ _1280_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6422_ _1854_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4517__B2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3634_ mod.registers.r10\[2\] _0602_ _0603_ mod.registers.r9\[2\] _0604_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _2707_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3565_ _3286_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ mod.registers.r1\[8\] _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6284_ _2944_ _2937_ _2945_ _2941_ _2742_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_fanout97_I net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3496_ _3177_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5235_ mod.des.des_dout\[22\] _2167_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3443__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__CLK net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _0727_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4983__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4117_ _1083_ _1084_ _1085_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5097_ mod.pc_2\[8\] _2042_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4048_ _1011_ _1012_ _1016_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_71_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4205__B1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ _2719_ _2721_ _2716_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__C2 mod.registers.r4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4851__S1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5181__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__B2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4449__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3798__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4747__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A3 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5743__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4787__C _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3350_ _3196_ _3197_ _3172_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4359__I _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _0886_ _0895_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _0069_ net113 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ mod.registers.r13\[10\] _2668_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4986__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ _2625_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4804_ _1659_ _1767_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4738__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4822__I _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5784_ mod.registers.r10\[7\] _2580_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4735_ _1437_ _1703_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3438__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4666_ _0802_ _1356_ _1364_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _1831_ _2856_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5163__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3617_ mod.registers.r9\[5\] _0427_ _0430_ mod.registers.r3\[5\] _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4597_ _0901_ _1565_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4910__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ _2978_ _2981_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3548_ _0441_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6267_ _2717_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _1786_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _2085_ _2876_ _2881_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5149_ _1932_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4977__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__CLK net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5154__A1 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3704__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__A1 mod.ldr_hzd\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3468__A1 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6406__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout147_I net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4196__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4520_ _1148_ _1149_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3943__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _0924_ _0790_ _0800_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3402_ mod.instr_2\[3\] _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4382_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _2816_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3333_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _2746_ mod.pc0\[12\] _2761_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _3155_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3721__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4959__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6954_ _0052_ net198 mod.ldr_hzd\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ _2399_ _2654_ _2660_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3631__A1 mod.registers.r6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _0386_ net172 mod.instr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__B2 mod.registers.r5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3596__C _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ _2556_ _2612_ _2616_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5384__A1 mod.registers.r2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4187__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5767_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4718_ _1343_ _1686_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_108_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ mod.registers.r8\[13\] _2522_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4649_ _1514_ _0945_ _1366_ _1477_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5687__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ _2961_ _2970_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4111__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5558__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__I _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5375__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5127__A1 mod.pc0\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3689__A1 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3541__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3861__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__B2 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6821__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5602__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3951_ _0724_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3613__A1 mod.registers.r11\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3613__B2 mod.registers.r2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4372__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6670_ _0174_ net98 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3882_ _0844_ _0845_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5621_ mod.registers.r7\[0\] _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4169__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6971__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _0717_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5118__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ _2254_ _2373_ _2376_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4434_ _1402_ _1403_ _1313_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4365_ _1333_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _1999_ _2766_ _2806_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3695__A4 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3316_ _3166_ _3168_ _3160_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_101_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1265_ _1070_ _0460_ _0452_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2746_ mod.pc0\[7\] _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3451__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3852__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3852__B2 mod.registers.r7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6397__A3 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__A1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6937_ _0035_ net195 mod.rd_3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5378__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6868_ _0369_ net191 mod.pc_1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ _2598_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _0303_ net110 mod.registers.r13\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3368__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3626__I _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3361__I _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6994__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5060__A3 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4859__B1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4323__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3531__B1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _1111_ _1112_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6076__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__I _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ mod.pc_2\[2\] _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4087__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_260 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_271 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_282 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_293 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _1627_ _1645_ _1385_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3598__B1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6722_ _0226_ net120 mod.registers.r8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3934_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A1 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3865_ mod.registers.r15\[10\] _0765_ _0766_ mod.registers.r12\[10\] _0835_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6653_ _0157_ net131 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5926__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ mod.registers.r6\[11\] _2460_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _0515_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6584_ _3139_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4562__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5535_ mod.registers.r5\[7\] _2405_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3365__A3 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5466_ mod.registers.r4\[3\] _2362_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3890__B _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4417_ _0949_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5397_ _2268_ _2315_ _2320_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6867__CLK net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4348_ _0828_ _0861_ _1253_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4277__I _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _1094_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4078__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _2736_ _1959_ _1965_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__B2 mod.registers.r10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5578__A1 mod.registers.r6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4250__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3761__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4069__A1 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4069__B2 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__A1 mod.registers.r13\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__B2 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__I _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6230__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5033__A3 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__B2 mod.registers.r7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3650_ _0595_ _0599_ _0613_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3694__C _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5741__A1 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3581_ _0530_ _0528_ _0539_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5320_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5251_ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ mod.registers.r3\[11\] _0694_ _0879_ mod.registers.r7\[11\] _1172_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3504__B1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5182_ _1907_ _2136_ _1377_ _0984_ _2072_ net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4133_ _1047_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ mod.registers.r11\[6\] _3202_ _3194_ mod.registers.r10\[6\] mod.registers.r2\[6\]
+ _3190_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout42_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _1388_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6705_ _0209_ net105 mod.registers.r7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3917_ _3172_ _3214_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4897_ mod.ldr_hzd\[15\] _1852_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3991__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6636_ _0140_ net78 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3848_ mod.registers.r4\[11\] _0419_ _3264_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3779_ _0747_ _0433_ _0661_ _0563_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6567_ _3118_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5518_ _2400_ _2389_ _2401_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6498_ _3087_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _2290_ _2349_ _2353_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3904__I _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout110 net112 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout121 net127 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout132 net133 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout154 net155 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout165 net166 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout176 net177 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout187 net188 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout198 net199 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5799__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__I0 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A1 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__B2 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5566__I _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__C _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6598__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3734__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5250__B _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout177_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4751_ _1228_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4765__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5962__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4380__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3702_ mod.registers.r6\[1\] _0503_ _0515_ mod.registers.r12\[1\] _0672_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4682_ _1444_ _1456_ _1151_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _3198_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6421_ _1813_ _3033_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5714__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3725__B1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6352_ _2985_ _2991_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3564_ _3282_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _2178_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6283_ mod.des.des_dout\[18\] _2900_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3724__I _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3495_ _3173_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _2181_ _1910_ _2174_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5165_ _2107_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ mod.registers.r15\[5\] _0485_ _3208_ mod.registers.r14\[5\] _1086_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5096_ mod.pc_2\[8\] _2042_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6905__CLK net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4047_ _0482_ _0483_ mod.registers.r1\[7\] _1014_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_72_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__B2 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5998_ mod.valid1 _2709_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5953__A1 mod.registers.r14\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ mod.pc_2\[1\] _1046_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6619_ _0123_ net84 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5705__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4692__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6197__A1 mod.pc_1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3809__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3707__B1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3544__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6121__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6928__CLK net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6970_ _0068_ net113 mod.registers.r15\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _2421_ _2667_ _2670_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4986__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6188__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5852_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4803_ _1769_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4199__B1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5935__A1 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _2546_ _2579_ _2583_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4734_ _1437_ _1703_ _1243_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4665_ _1406_ _1362_ _1533_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6404_ _0687_ _2956_ _3024_ _2855_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3616_ mod.registers.r15\[5\] _0434_ _0436_ mod.registers.r12\[5\] _0586_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5163__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__A1 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _1541_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6335_ _0636_ _2975_ _2979_ mod.instr\[12\] _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_1_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3547_ _0439_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4910__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6112__A1 _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ mod.instr\[14\] _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3478_ _0444_ _0445_ _0410_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5217_ _1786_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4674__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6197_ mod.pc_1\[10\] _2877_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _1907_ _2090_ _2105_ _3156_ _2106_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_96_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5079_ _1896_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6351__A1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3364__I _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__B1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4665__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3468__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6406__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4968__A2 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5090__B2 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5754__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3943__A3 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4450_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6750__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3401_ _3252_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4381_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6120_ _1925_ _2048_ _2051_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3332_ _3181_ _3167_ _3183_ _3184_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2722_ _2114_ _2117_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _1385_ _1621_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_22_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _0051_ net198 mod.ldr_hzd\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4959__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5904_ mod.registers.r13\[3\] _2656_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6884_ _0385_ net172 mod.instr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5835_ mod.registers.r11\[10\] _2613_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5908__A1 mod.registers.r13\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3449__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5766_ _2570_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4989__B _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4592__B1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _0497_ _0827_ _0841_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5664__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5697_ _2431_ _2521_ _2523_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4648_ _1095_ _1370_ _1548_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6333__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__B2 mod.instr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4895__A1 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ mod.instr_2\[6\] _2968_ _2963_ mod.instr\[6\] _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _2918_ _2913_ _2919_ _2917_ _2911_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4647__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3912__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5574__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3689__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A1 mod.instr_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4918__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4638__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3861__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5749__I _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A1 mod.pc_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _3248_ _0916_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3613__A2 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3881_ _0777_ _0847_ _0849_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_32_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5620_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4023__C1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4169__A3 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5551_ _2267_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _1467_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5482_ mod.registers.r4\[9\] _2374_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4433_ _0525_ _0461_ _0592_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4341__A3 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4364_ _1205_ _0799_ _3262_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6103_ _2767_ _2805_ _2778_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3315_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4295_ _0578_ _0494_ _1069_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_86_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _2736_ _2032_ _2035_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout72_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6646__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5054__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5659__I _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _0034_ net184 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4801__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3604__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6796__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6867_ _0368_ net193 mod.pc_1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ _2538_ _2599_ _2605_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5357__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6798_ _0302_ net113 mod.registers.r13\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3368__A1 mod.registers.r14\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3368__B2 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5749_ _2275_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3907__A3 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5109__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A1 mod.registers.r1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6545__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4020__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4859__B2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3531__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3531__B2 mod.registers.r10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ _1033_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_250 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_261 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_272 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_283 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_294 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5036__A1 mod.pc0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4244__C1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0699_ _0710_ _3223_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3598__A1 mod.registers.r10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6721_ _0225_ net105 mod.registers.r8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3598__B2 mod.registers.r2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3933_ _3230_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6652_ _0156_ net83 mod.registers.r3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5339__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3864_ mod.registers.r9\[10\] _0751_ _0752_ mod.registers.r3\[10\] _0834_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6536__A1 mod.registers.r15\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _2425_ _2459_ _2463_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6583_ net17 mod.des.des_dout\[27\] _3137_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _0514_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3727__I _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5534_ _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3770__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5465_ _2194_ _2360_ _2365_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4416_ _0943_ _1380_ _1381_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ mod.registers.r2\[11\] _2316_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4347_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4278_ _1033_ _1049_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4078__A2 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2728_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5027__A1 mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3589__A1 mod.registers.r14\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _0017_ net183 mod.pc_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3589__B2 mod.registers.r6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4250__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6527__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3637__I _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3761__A1 mod.registers.r8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3761__B2 mod.registers.r10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5852__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6550__I1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3372__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5266__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4069__A2 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3816__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3547__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout122_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3580_ _0540_ _0543_ _0546_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ mod.des.des_dout\[24\] _2167_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _1168_ _1169_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3504__A1 mod.registers.r8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5181_ _1907_ _2136_ _1435_ _1001_ _2072_ net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4132_ _1050_ _1073_ _1096_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_96_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__A1 mod.des.des_dout\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4063_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4480__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _1932_ _1604_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6704_ _0208_ net59 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3916_ _0880_ _0881_ _0883_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4896_ _1848_ _1860_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6635_ _0139_ net78 mod.registers.r2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3991__B2 mod.registers.r2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3847_ mod.registers.r11\[11\] _0505_ _0412_ mod.registers.r2\[11\] _0817_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6834__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6566_ _3128_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3778_ mod.registers.r15\[12\] _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4535__A3 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3743__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5517_ mod.registers.r5\[3\] _2391_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6497_ mod.des.des_dout\[9\] net7 _3085_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5448_ mod.registers.r3\[14\] _2350_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5496__A1 mod.registers.r4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6984__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout100 net102 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5379_ _2303_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout111 net112 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout122 net124 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout133 net150 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout144 net148 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout155 net160 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout166 net167 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout177 net178 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout188 net194 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__I1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4471__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6008__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5971__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3982__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3734__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3734__B2 mod.registers.r9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4926__I _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5757__I _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ _1247_ _1706_ _1707_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3701_ mod.registers.r13\[1\] _0520_ _3272_ mod.registers.r8\[1\] _0671_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4681_ _1279_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6420_ _3034_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3632_ _3194_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6351_ mod.funct7\[0\] _2989_ _2986_ mod.instr\[18\] _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3725__B2 mod.registers.r7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3563_ mod.registers.r8\[7\] _0531_ _0532_ mod.registers.r10\[7\] _0533_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5302_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6282_ mod.instr\[18\] _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3494_ _3265_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3740__A4 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5233_ mod.pc_2\[1\] _2182_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5164_ _1727_ _1737_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4115_ mod.registers.r8\[5\] _3204_ _3198_ mod.registers.r9\[5\] _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _1970_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ mod.registers.r3\[7\] _1013_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4453__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3896__B _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5997_ _2712_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4948_ _1206_ _3259_ _1077_ _3263_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4504__C _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4879_ _0490_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6618_ _0122_ net85 mod.registers.r1\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6549_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5181__A3 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__I _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A3 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4444__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5641__A1 mod.registers.r7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__I _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A1 mod.registers.r5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3707__B2 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6201__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A1 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3560__I mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4435__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5920_ mod.registers.r13\[9\] _2668_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5851_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4802_ _1182_ _1397_ _1641_ _1330_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4199__A1 mod.registers.r11\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4199__B2 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5782_ mod.registers.r10\[6\] _2580_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4733_ _1442_ _1682_ _1675_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5148__B1 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _1541_ _1612_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5699__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ mod.ri_3 _2867_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3615_ _0581_ _0582_ _0583_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4595_ _1357_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3735__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6334_ _2978_ _2980_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3546_ mod.registers.r15\[6\] _0514_ _0515_ mod.registers.r12\[6\] _0516_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4910__A3 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6265_ _2930_ _2925_ _2931_ _2929_ _2923_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3477_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5950__I _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4123__A1 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6196_ _2872_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5871__A1 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4674__A2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _1171_ _1176_ _1929_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3470__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _1909_ _1511_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5623__A1 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ mod.registers.r3\[14\] _0959_ _0960_ mod.registers.r2\[14\] _0999_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3634__B1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4114__A1 mod.registers.r4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__B2 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3380__I _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5614__A1 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__B _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3555__I _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4353__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3400_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout202_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ _0621_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3331_ mod.instr_2\[14\] _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _2759_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _1949_ _1967_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3864__B1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _0050_ net174 mod.ldr_hzd\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3616__B1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5081__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _2396_ _2654_ _2659_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6883_ _0384_ net171 mod.instr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5834_ _2554_ _2612_ _2615_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5765_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4716_ _1317_ _1409_ _1592_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5696_ mod.registers.r8\[12\] _2522_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _1074_ _1337_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3465__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4578_ _0930_ _0932_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _2961_ _2969_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3529_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ mod.des.des_dout\[9\] _2909_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5844__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6179_ _2860_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3855__B1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6021__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__CLK net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4583__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5076__B _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3375__I mod.funct3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A2 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6088__A1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5835__A1 mod.registers.r11\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__B1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3310__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6260__A1 mod.des.des_dout\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5063__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout152_I net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3880_ _0846_ _0632_ mod.registers.r8\[8\] _0638_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4023__B1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__C2 mod.registers.r10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _2425_ _2418_ _2426_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4501_ _0925_ _1410_ _1414_ _1469_ _1470_ _1315_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_117_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5481_ _2245_ _2373_ _2375_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4432_ _1401_ _1310_ _0576_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4363_ _0692_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A1 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6102_ _2801_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3314_ mod.instr_2\[16\] _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _0625_ _0680_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5826__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4629__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _2743_ _2748_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5005__I mod.pc_2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout65_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0033_ net185 mod.ri_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6866_ _0367_ net189 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ mod.registers.r11\[3\] _2601_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _0301_ net109 mod.registers.r13\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5675__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3368__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _2558_ _2551_ _2559_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _2408_ _2509_ _2512_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4317__A1 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3923__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3540__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5817__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3828__B1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6740__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4308__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3531__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_240 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6365__B _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_251 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_262 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3834__A3 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_273 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_284 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_295 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6084__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6233__B2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _1931_ _1948_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4244__B1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4244__C2 mod.registers.r15\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4795__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3932_ _0457_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6720_ _0224_ net60 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3598__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _0155_ net80 mod.registers.r3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3863_ _0829_ _0830_ _0831_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6536__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5602_ mod.registers.r6\[10\] _2460_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6582_ _3138_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3794_ _0760_ _0761_ _0762_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5533_ _2235_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3770__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5464_ mod.registers.r4\[2\] _2362_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4415_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5395_ _2261_ _2315_ _2319_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4346_ _0801_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6472__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _2733_ _2735_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6763__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3589__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _0016_ net169 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6849_ _0350_ net158 mod.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3761__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__C1 mod.registers.r11\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4433__B _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout115_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4200_ mod.registers.r6\[11\] _0700_ _0889_ mod.registers.r13\[11\] _1170_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3504__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _2107_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4131_ _1097_ _1049_ _1098_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A2 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4062_ _1030_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6206__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _1385_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _0207_ net100 mod.registers.r7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3915_ mod.registers.r15\[4\] _0884_ _0600_ mod.registers.r6\[4\] _0603_ mod.registers.r9\[4\]
+ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_4895_ _1861_ _1863_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ _0138_ net86 mod.registers.r2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3991__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3846_ mod.registers.r14\[11\] _0502_ _0503_ mod.registers.r6\[11\] _0816_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6565_ mod.des.des_dout\[20\] net5 _3124_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3777_ mod.registers.r12\[12\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3743__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ _2399_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6496_ _3086_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5447_ _2284_ _2349_ _2352_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5496__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5378_ _2301_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout101 net102 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout112 net118 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4329_ _0991_ _1296_ _1297_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout134 net137 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout145 net147 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout156 net159 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout167 net168 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout178 net179 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout189 net193 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4846__I2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3734__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3558__I _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ mod.registers.r1\[1\] _0521_ _0412_ mod.registers.r2\[1\] _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4680_ _1648_ _1649_ _1128_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3631_ mod.registers.r6\[2\] _0600_ _3189_ mod.registers.r5\[2\] mod.registers.r2\[2\]
+ _3191_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6350_ _2985_ _2990_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3725__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3562_ _3278_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ mod.des.des_dout\[29\] _2188_ _2240_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ _2942_ _2937_ _2943_ _2941_ _2935_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3493_ _0454_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5232_ _1793_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3489__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _1196_ _1199_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A1 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4114_ mod.registers.r4\[5\] _0465_ _3194_ mod.registers.r10\[5\] _1084_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5094_ _1909_ _1674_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4338__B _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4045_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _1789_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4878_ mod.instr_2\[6\] _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6617_ _0121_ net84 mod.registers.r1\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6951__CLK net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ _0791_ _0796_ _0797_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_20_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3716__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ mod.des.des_counter\[2\] _1906_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_106_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6479_ mod.des.des_dout\[1\] net17 _3075_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4141__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__A1 mod.instr_2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3378__I mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6354__B1 _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3707__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__I _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4132__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout182_I net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__B _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5850_ _2357_ _2624_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _1180_ _1670_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6974__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4199__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5781_ _2544_ _2579_ _2582_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4732_ _1256_ _1678_ _1700_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5148__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ _0989_ _1538_ _1345_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4621__B _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5699__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3614_ mod.registers.r4\[5\] _0418_ _3236_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6402_ _3021_ _3022_ _3023_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4594_ _0989_ _1316_ _1341_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3545_ _0436_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6333_ _1808_ _2975_ _2979_ mod.instr\[11\] _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4910__A4 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__I1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6264_ mod.des.des_dout\[13\] _2921_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3476_ _0444_ _0445_ _3281_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_89_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4123__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _2066_ _2876_ _2879_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5871__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5146_ _2101_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3882__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _2037_ _2038_ _2039_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4028_ mod.registers.r15\[14\] _0964_ _0968_ mod.registers.r8\[14\] _0998_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3634__A1 mod.registers.r10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3634__B2 mod.registers.r9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ net11 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6503__S _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4898__C2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3570__B1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5311__A1 mod.des.des_dout\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4114__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6847__CLK net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A3 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6997__CLK net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3928__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4050__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6212__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4889__B1 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4353__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4105__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3571__I _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _3225_ _1950_ _1966_ _1904_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__B2 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _0049_ net175 mod.ldr_hzd\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5498__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3616__A1 mod.registers.r15\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5902_ mod.registers.r13\[2\] _2656_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6882_ _0383_ net178 mod.instr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ mod.registers.r11\[9\] _2613_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6318__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4715_ _1436_ _1680_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3746__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5695_ _2503_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__I _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4646_ _1518_ _1269_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_163_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5541__A1 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _1076_ _1099_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3552__B1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _2967_ _2968_ _2963_ mod.instr\[5\] _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3528_ _0457_ _3257_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6247_ mod.instr\[9\] _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3459_ _3289_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__C1 _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3855__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6178_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3855__B2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5129_ _3225_ _2074_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6021__A2 mod.pc0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4032__A1 mod.funct7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__B1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5780__A1 mod.registers.r10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__B1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5532__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3543__B1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5092__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3605__B _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4638__A3 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5835__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3846__A1 mod.registers.r14\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__B2 mod.registers.r6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5599__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6207__I mod.instr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A2 _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout145_I net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__A1 mod.registers.r4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4023__B2 mod.registers.r1\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _1403_ _1413_ _0496_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5480_ mod.registers.r4\[8\] _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _0667_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5523__A1 mod.registers.r5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__B1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4362_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__I _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ _1998_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3313_ _3161_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4293_ _1260_ _1261_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _2746_ mod.pc0\[6\] _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6117__I _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6934_ _0032_ net184 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4262__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6865_ _0366_ net190 mod.pc_1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5816_ _2536_ _2599_ _2604_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6796_ _0300_ net44 mod.registers.r12\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5762__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5747_ mod.registers.r9\[11\] _2552_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6692__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ mod.registers.r8\[5\] _2510_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5514__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0576_ _0592_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3828__A1 mod.registers.r8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3828__B2 mod.registers.r15\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5753__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3386__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3764__B1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5505__A1 mod.registers.r5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4010__I _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4945__I _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_230 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_241 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_252 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_263 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_274 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_285 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A2 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_296 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4244__A1 mod.registers.r3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _3225_ _1933_ _1947_ _1904_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4244__B2 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5776__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6650_ _0154_ net83 mod.registers.r3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ mod.registers.r4\[10\] _0420_ _3265_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5601_ _2422_ _2459_ _2462_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5744__A1 mod.registers.r9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ net16 mod.des.des_dout\[26\] _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3793_ mod.registers.r4\[13\] _0738_ _3238_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5532_ _2411_ _2404_ _2412_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ _2186_ _2360_ _2364_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5394_ mod.registers.r2\[10\] _2316_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0809_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4276_ _0940_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6908__CLK net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2734_ mod.pc0\[2\] _2731_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _0015_ net169 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4786__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _0349_ net157 mod.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4538__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _0283_ net81 mod.registers.r11\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3934__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4171__B1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__C2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3521__I0 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6215__A2 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4005__I _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__B1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3844__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6220__I _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__A1 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4701__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4130_ _1076_ _1099_ _1075_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ _1029_ _1022_ _1026_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_56_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A3 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6206__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4217__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5965__A1 mod.registers.r14\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _0599_ _0613_ _3223_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _0206_ net100 mod.registers.r7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3914_ _0485_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4894_ mod.ldr_hzd\[6\] _1858_ _1854_ mod.ldr_hzd\[5\] _1851_ mod.ldr_hzd\[7\] _1864_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_20_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _0137_ net77 mod.registers.r2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5717__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3845_ mod.registers.r8\[11\] _0531_ _0500_ mod.registers.r10\[11\] _0815_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3728__B1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _3127_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3776_ _0521_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5515_ _2198_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6495_ mod.des.des_dout\[8\] net6 _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3754__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ mod.registers.r3\[13\] _2350_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6730__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _2199_ _2302_ _2308_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout102 net108 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout113 net117 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3900__B1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout135 net137 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4328_ _1296_ _1297_ _0992_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout146 net148 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout157 net159 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3703__B _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout168 net181 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout179 net180 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4259_ _1226_ _1201_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6880__CLK net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4456__B2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__I3 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4208__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4759__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5956__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 mod.pc_1\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6040__I _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4696__S _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3742__I0 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 mod.registers.r14\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3839__I _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3630_ _3185_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6372__A1 mod.pc_1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6753__CLK net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3574__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3561_ _3271_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _2213_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6124__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ mod.des.des_dout\[17\] _2933_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3492_ _0461_ _0453_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5231_ _1793_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4686__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3489__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ _2109_ _2119_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4150__A3 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__B _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ mod.registers.r12\[5\] _0887_ _3185_ mod.registers.r6\[5\] _1083_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5093_ _1908_ _2040_ _2053_ _0001_ _2054_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_96_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4044_ _3166_ _3216_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout40_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__I _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1789_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _1838_ _1841_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _0120_ net89 mod.registers.r1\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ mod.registers.r8\[15\] _0729_ _0765_ mod.registers.r15\[15\] _0798_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6363__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _2441_ _3112_ _3117_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3759_ _3272_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4913__A2 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _3076_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _2229_ _2337_ _2341_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__B _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__I _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6626__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__A2 mod.instr_2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5874__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6354__A1 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3394__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__B2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__B _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__B2 _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout175_I net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _1181_ _1484_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ mod.registers.r10\[5\] _2580_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4731_ _1700_ _1256_ _1678_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ _0925_ _1561_ _1630_ _1306_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__5148__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _2715_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3613_ mod.registers.r11\[5\] _3291_ _0411_ mod.registers.r2\[5\] _0583_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4593_ _1559_ _1562_ _1327_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _2950_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3544_ _0434_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6263_ mod.instr\[13\] _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3475_ _0426_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5214_ _2142_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6194_ mod.pc_1\[9\] _2877_ _2873_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ mod.pc0\[11\] _1892_ _1901_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3882__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _1008_ _1020_ _1985_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5959__I _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4027_ mod.registers.r6\[14\] _0966_ _0967_ mod.registers.r5\[14\] _0997_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3634__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4831__A1 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3479__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _2441_ _2700_ _2705_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4434__I1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _1884_ _1889_ _1895_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5694__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5139__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3570__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3570__B2 mod.registers.r12\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__B _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3389__I _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__C1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A1 mod.pc_2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6941__CLK net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6950_ _0048_ net174 mod.ldr_hzd\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3616__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5901_ _2393_ _2654_ _2658_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6881_ _0382_ net178 mod.instr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5832_ _2550_ _2612_ _2614_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _2299_ _2499_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4632__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4714_ _1243_ _1683_ _1433_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6318__A1 mod.instr_2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _2501_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ _1518_ _1514_ _1241_ _0940_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5019__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3927__I0 mod.funct7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _1306_ _1544_ _1545_ _1309_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5541__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3552__A1 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _2955_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3552__B2 mod.registers.r1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3762__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6246_ _2915_ _2913_ _2916_ _2917_ _2911_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3458_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4501__B1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4501__C2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6177_ _2857_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3389_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3855__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _2084_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5059_ _1037_ _1042_ _1985_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6313__I _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6309__A1 mod.instr_2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A1 mod.registers.r14\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3791__B2 mod.registers.r6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5532__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3543__A1 mod.registers.r9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4768__I _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__I0 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3543__B2 mod.registers.r3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6964__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A1 mod.pc_2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3846__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5048__A1 mod.pc_2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4008__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__A1 mod.ins_ldr_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6223__I _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout138_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _0726_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A1 mod.registers.r14\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__B _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4678__I _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__B2 mod.registers.r6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _0917_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3582__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6100_ _2802_ _2769_ mod.pc\[5\] _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3312_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4292_ _0723_ _0666_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _2736_ _2016_ _2019_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5302__I _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6933_ _0031_ net184 mod.valid_out3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4262__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6864_ _0365_ net190 mod.pc_1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5815_ mod.registers.r11\[2\] _2601_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3757__I mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ _0299_ net81 mod.registers.r12\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__CLK net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _2267_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5762__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5677_ _2403_ _2509_ _2511_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4628_ _1313_ _0555_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _1320_ _1354_ _1344_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5278__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6229_ _2891_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3828__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6308__I _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4253__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5202__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3764__A1 mod.registers.r14\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3764__B2 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6199__B _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4498__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3516__A1 mod.registers.r15\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_220 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_231 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_242 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6218__I _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_253 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_264 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_275 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_286 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_297 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _0878_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__B _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ mod.registers.r11\[10\] _3292_ _0413_ mod.registers.r2\[10\] _0831_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3577__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ mod.registers.r6\[9\] _2460_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6580_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3792_ mod.registers.r11\[13\] _0735_ _0736_ mod.registers.r2\[13\] _0762_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5744__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ mod.registers.r5\[6\] _2405_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ mod.registers.r4\[1\] _2362_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4413_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5393_ _2254_ _2315_ _2318_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4180__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ _1309_ _1312_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6457__B1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4275_ _1240_ _1243_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6014_ _2728_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout70_I net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A1 mod.registers.r8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6916_ _0014_ net169 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _0348_ net153 mod.pc0\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _0282_ net77 mod.registers.r11\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5729_ _2228_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4171__B2 mod.registers.r5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4474__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3521__I1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3682__B1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3737__A1 mod.registers.r11\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3737__B2 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__A1 mod.registers.r10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4956__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4060_ _1022_ _1026_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6682__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4870__C1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5787__I _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5414__A1 mod.registers.r3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _1908_ _1910_ _1928_ _0001_ _1930_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__5965__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3976__A1 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _0205_ net59 mod.registers.r7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3913_ mod.registers.r5\[4\] _0882_ _0706_ mod.registers.r8\[4\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4893_ mod.ldr_hzd\[4\] _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6632_ _0136_ net87 mod.registers.r2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3844_ _0557_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3728__A1 mod.registers.r4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ mod.des.des_dout\[19\] net4 _3124_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3728__B2 mod.registers.r1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3775_ _0520_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6390__A2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _2397_ _2389_ _2398_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6494_ _3074_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5445_ _2276_ _2349_ _2351_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4153__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ mod.registers.r2\[3\] _2304_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout103 net107 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3900__A1 mod.registers.r9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _1003_ _1232_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout114 net117 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3900__B2 mod.registers.r3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout125 net127 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout136 net137 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout147 net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout158 net159 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _1221_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout169 net173 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4456__A2 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5653__A1 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ mod.registers.r14\[10\] _0891_ _0703_ mod.registers.r9\[10\] mod.registers.r2\[10\]
+ _0893_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4534__C _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4759__A3 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4106__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3719__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__I _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6908__D _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3742__I1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4447__A2 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4383__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout218_I net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3560_ mod.pc_2\[7\] _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4135__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _2164_ _2177_ _2180_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6387__B _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__B _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _1985_ _1218_ _2118_ _1969_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__B1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ _1079_ _1080_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_68_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ _1131_ _1142_ _1929_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A1 mod.registers.r7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _3209_ _3217_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ mod.valid0 _2709_ _2151_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_52_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4945_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4071__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _1842_ _1843_ _1844_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_20_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3827_ mod.registers.r11\[15\] _0735_ _0738_ mod.registers.r4\[15\] _0736_ mod.registers.r2\[15\]
+ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6615_ _0119_ net90 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3765__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6546_ mod.registers.r15\[15\] _3113_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3758_ _3266_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6477_ mod.des.des_dout\[0\] net16 _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5980__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3689_ mod.registers.r9\[3\] _0544_ _0545_ mod.registers.r3\[3\] _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4126__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ mod.registers.r3\[6\] _2338_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ mod.des.des_dout\[36\] _2220_ _2292_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_87_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3885__B1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5929__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6051__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 mod.registers.r12\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3624__B _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3628__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5093__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__B2 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4455__B _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout168_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _1437_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__B1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _1318_ _1321_ _0626_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6400_ _1886_ _1798_ _3249_ _2858_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6870__CLK net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3612_ mod.registers.r14\[5\] _3282_ _3286_ mod.registers.r6\[5\] _0582_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _0692_ _1560_ _1561_ _0626_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6331_ _2759_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3543_ mod.registers.r9\[6\] _0511_ _0512_ mod.registers.r3\[6\] _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6262_ _2927_ _2925_ _2928_ _2929_ _2923_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3474_ _0425_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5856__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _2050_ _2876_ _2878_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3867__B1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5144_ _2102_ _2041_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 mod.registers.r6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3882__A3 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _1987_ _2024_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__B1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _0993_ _0994_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5040__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5977_ mod.registers.r14\[15\] _2701_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3398__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _1893_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _0640_ _1816_ _1821_ _0848_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _3094_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3570__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 mod.registers.r11\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5215__I _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5075__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__B1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4035__C2 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6893__CLK net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4050__A3 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4889__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5838__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4105__A4 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__I mod.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4964__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5900_ mod.registers.r13\[1\] _2656_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6880_ _0381_ net176 mod.instr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6015__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ mod.registers.r11\[8\] _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5762_ _2568_ _2561_ _2569_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4041__A3 mod.registers.r8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4713_ _1442_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6318__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5693_ _2428_ _2515_ _2520_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _1609_ _1610_ _1612_ _1566_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3927__I1 mod.funct7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4575_ _1468_ _1501_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6314_ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3526_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3552__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _2891_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3457_ _0424_ _3269_ _0425_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6176_ _1962_ _2859_ _2866_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3388_ _3227_ _3229_ _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ mod.pc0\[10\] _1922_ _1923_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_29_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__A2 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ _1987_ _2007_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input13_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4804__A2 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4009_ mod.registers.r14\[15\] _0977_ _0978_ mod.registers.r7\[15\] _0979_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A3 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3791__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3953__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4591__I1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3543__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5296__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5048__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4733__B _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6639__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _1328_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3534__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6789__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3311_ _3160_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _0807_ _0650_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _2722_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5287__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6932_ _0030_ net182 mod.pc_2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _0364_ net191 mod.pc_1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5814_ _2534_ _2599_ _2603_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6794_ _0298_ net79 mod.registers.r12\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__A2 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5745_ _2556_ _2551_ _2557_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4970__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5676_ mod.registers.r8\[4\] _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4627_ _0593_ _0860_ _0875_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3773__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__C1 mod.registers.r3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4558_ _1318_ _1321_ _1406_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3509_ mod.registers.r12\[1\] _0476_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4489_ _1228_ _1222_ _1458_ _1285_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6228_ mod.des.des_dout\[4\] _2896_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _2850_ _2852_ _2818_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4789__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5450__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3948__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5202__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3764__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6931__CLK net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3516__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6466__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_221 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_232 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_243 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_254 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_265 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_276 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4019__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_287 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_298 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3858__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3452__A1 mod.registers.r4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout150_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ mod.registers.r14\[10\] _0732_ _0733_ mod.registers.r6\[10\] _0830_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3791_ mod.registers.r14\[13\] _3283_ _3287_ mod.registers.r6\[13\] _0761_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5461_ _2177_ _2360_ _2363_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4412_ _0942_ _0932_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3507__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5392_ mod.registers.r2\[9\] _2316_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ _0923_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4180__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__B2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4274_ _1239_ _1004_ _1238_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _2726_ _1947_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout63_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _0013_ net144 mod.instr_2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3768__I _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6846_ _0347_ net153 mod.pc0\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6954__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _0281_ net77 mod.registers.r11\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3989_ _3165_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5728_ _2544_ _2541_ _2545_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5659_ _2149_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4171__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3452__B _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3682__A1 mod.registers.r8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3682__B2 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4162__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4458__B _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6229__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6827__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout198_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3673__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__C2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__B _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _0470_ _0488_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6700_ _0204_ net39 mod.registers.r6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3912_ _3188_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3976__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4892_ _1856_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _0135_ net88 mod.registers.r2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5178__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3843_ _0556_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3728__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6562_ _3126_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3774_ mod.registers.r7\[12\] _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5513_ mod.registers.r5\[2\] _2391_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6493_ _3084_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ mod.registers.r3\[12\] _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5350__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _2194_ _2302_ _2307_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout104 net107 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4326_ _1287_ _1295_ _1236_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3900__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout115 net117 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout126 net127 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout137 net141 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__A1 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout148 net149 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4257_ _1226_ _1201_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout159 net160 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_68_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5653__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4188_ mod.registers.r6\[10\] _0700_ _0705_ mod.registers.r11\[10\] _1158_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5405__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3498__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6829_ _0000_ _0004_ net206 mod.des.des_counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3719__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5218__I _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4144__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3352__B1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6049__I _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4907__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4383__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__A1 mod.registers.r6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout113_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3490_ _0455_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4135__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _2114_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__A1 mod.registers.r14\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3894__B2 mod.registers.r6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ mod.registers.r5\[5\] _3188_ _3211_ mod.registers.r13\[5\] _1081_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5091_ _2049_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _0951_ _3216_ mod.registers.r4\[7\] _1010_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5635__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7005__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5993_ _2710_ _2714_ _2716_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1911_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4071__A1 mod.registers.r12\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__B2 mod.registers.r13\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4875_ _1802_ _1834_ _1835_ _1810_ _1836_ _1804_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__6422__I _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _0118_ net90 mod.registers.r1\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3826_ _0792_ _0793_ _0794_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _2438_ _3112_ _3116_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5571__A1 mod.registers.r5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ mod.pc_2\[12\] _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _3074_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3688_ mod.registers.r7\[3\] _0548_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ _2218_ _2337_ _2340_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5323__A1 mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3781__I _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5358_ _2226_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3885__A1 mod.registers.r14\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3885__B2 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ _0873_ _1124_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5289_ _1935_ _2208_ _2226_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6051__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4062__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3956__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6332__I _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4365__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3691__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4668__A3 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__A2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3628__A1 mod.registers.r4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6290__A2 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6507__I _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5411__I _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3643__A4 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A1 mod.registers.r5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__B2 mod.registers.r7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _1628_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3611_ mod.registers.r8\[5\] _3271_ _3278_ mod.registers.r10\[5\] _0581_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4356__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__A1 mod.registers.r5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4591_ _0666_ _1251_ _0667_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6330_ _2971_ _2977_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3542_ _0430_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6398__B _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4108__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ net13 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3473_ mod.registers.r5\[0\] _0440_ _0442_ mod.registers.r7\[0\] _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5856__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5212_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3867__A1 mod.registers.r13\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6192_ mod.pc_1\[8\] _2877_ _2873_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3867__B2 mod.registers.r1\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5143_ mod.pc\[11\] _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ _1969_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3619__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3619__B2 mod.registers.r1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__A2 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4025_ mod.registers.r11\[14\] _0974_ _0980_ mod.registers.r13\[14\] _0995_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4292__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _2438_ _2700_ _2704_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4044__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3776__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _1823_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6592__I0 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4789_ _1281_ _1650_ _1741_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6528_ _3092_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _1802_ _3058_ _3059_ _3044_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5231__I _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A1 mod.registers.r15\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4035__B2 mod.registers.r6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5783__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4586__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 mod.registers.r5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__I0 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__B1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6011__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__A2 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6237__I _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout180_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__A2 mod.pc0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _2600_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ mod.registers.r9\[15\] _2562_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4577__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A1 mod.registers.r10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _1518_ _1096_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4041__A4 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5692_ mod.registers.r8\[11\] _2516_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4329__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _1501_ _1419_ _0776_ _0803_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6574__I0 mod.des.des_dout\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3537__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ _1312_ _1319_ _0593_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1861_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3525_ _0464_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ mod.des.des_dout\[8\] _2909_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3456_ mod.instr_2\[10\] _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3387_ _3233_ _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ mod.pc_1\[3\] _2861_ _2864_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _2085_ _1897_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4376__B _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _1969_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4265__A1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _3170_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _2680_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A1 mod.registers.r5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4740__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__I _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6710__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3700__B1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6057__I _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6860__CLK net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5756__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4559__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3767__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6181__A1 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__I mod.pc_2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3310_ _3161_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4290_ _1062_ _1063_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4196__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6931_ _0029_ net182 mod.pc_2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4798__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _0363_ net189 mod.pc_1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ mod.registers.r11\[1\] _2601_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5747__A1 mod.registers.r9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6793_ _0297_ net79 mod.registers.r12\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4215__I _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5744_ mod.registers.r9\[10\] _2552_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4970__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5675_ _2503_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _1327_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6733__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4183__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4183__C2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ _1524_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3508_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4488_ _1444_ _1456_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6227_ mod.instr\[4\] _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3439_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4486__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6883__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _2850_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5109_ _1109_ _1120_ _1929_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6089_ _2783_ _2785_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4238__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5738__A1 mod.registers.r9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4410__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__I _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A1 mod.registers.r13\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput30 net30 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_222 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_233 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_244 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_255 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_266 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_277 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_288 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_299 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5977__A1 mod.registers.r14\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6606__CLK net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3452__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout143_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3790_ mod.registers.r8\[13\] _3273_ _3279_ mod.registers.r10\[13\] _0760_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6756__CLK net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6250__I mod.instr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ mod.registers.r4\[0\] _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0943_ _1377_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5901__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2245_ _2315_ _2317_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4342_ _0527_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4919__B mod.valid0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4273_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6012_ _2730_ _1928_ _2732_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

